** sch_path: /home/gmaranhao/pdk/IHP-Open-PDK/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/sp_mim_cap.sch
**.subckt sp_mim_cap
R1 in GND 1Meg m=1
V1 in GND dc 0 ac 1 portnum 1 z0 50
R2 out GND 1Meg m=1
V2 out GND dc 0 ac 0 portnum 2 z0 50
XC1 out in cap_cmim W=7.0e-6 L=7.0e-6 MF=1
**** begin user architecture code


.control
save all
sp lin 500 1e9 100e9 0
let Cseries = 1e+15/(2*PI*frequency*imag(1/Y_2_1))
let Rseries = -real(1/Y_2_1)
write sp_mim_cap.raw
.endc



.lib /home/gmaranhao/pdk/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ

**** end user architecture code
**.ends
.GLOBAL GND
.end
