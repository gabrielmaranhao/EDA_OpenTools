** sch_path: /home/gmaranhao/Desktop/ihp130_work/nmos_idvd.sch
**.subckt nmos_idvd
Vds vd GND 0
V3 net2 GND 0
Vs net1 GND 0
Vgb vg GND 700m
XM1 vd vg net1 net2 sg13_lv_nmos W=10.0u L=0.12u ng=1 m=1
**** begin user architecture code



.control
pre_osdi ./psp103_nqs.osdi
save all

dc Vds 0.001 1.5 1m

let gmd = deriv(i(Vs))
save gmd

write nmos_idvd.raw

.endc




.lib /home/gmaranhao/pdk/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
