* NGSPICE file created from bias.ext - technology: sky130A

.subckt bias IREF AVDD AVSS VB3 VB4 VB2 VB1
X0 a_9838_205# VB2.t45 VB4.t10 AVSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1 AVSS.t179 AVSS.t177 AVSS.t178 AVSS.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2 a_8132_2488# IREF.t10 VB1.t0 AVSS.t194 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3 a_4970_1009# VB1.t65 VB1.t66 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X4 a_9838_2488# IREF.t11 VB1.t4 AVSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X5 a_10519_5228# VB4.t15 AVDD.t7 AVDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X6 AVSS.t176 AVSS.t174 AVSS.t175 AVSS.t33 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X7 AVSS.t173 AVSS.t170 AVSS.t172 AVSS.t171 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X8 AVSS.t169 AVSS.t168 AVSS.t169 AVSS.t59 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X9 a_8132_1583# IREF.t4 IREF.t5 AVSS.t194 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X10 a_2712_n77# VB1.t75 VB2.t9 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X11 AVDD.t126 VB1.t76 a_3744_4980# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X12 a_9838_1583# IREF.t8 IREF.t9 AVSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X13 VB4.t9 VB4.t8 a_10777_6298# AVDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X14 a_2712_4093# VB1.t77 VB2.t0 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X15 AVDD.t420 AVDD.t419 AVDD.t420 AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X16 a_2002_6484# VB1.t78 VB2.t31 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X17 AVDD.t125 VB1.t79 a_3744_2103# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X18 AVDD.t124 VB1.t80 a_2002_5597# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X19 AVDD.t123 VB1.t81 a_2712_5597# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X20 a_4970_n77# VB1.t82 VB3.t27 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X21 a_3744_4980# VB1.t83 VB3.t4 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X22 AVDD.t122 VB1.t84 a_4970_1009# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X23 a_10777_6298# VB4.t16 a_10519_6298# AVDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X24 a_4970_n2468# VB1.t85 VB2.t7 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X25 AVDD.t121 VB1.t86 a_4970_n3085# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X26 VB2.t28 VB1.t87 a_1486_6484# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X27 a_3744_2103# VB1.t5 VB1.t6 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X28 VB2.t34 VB1.t88 a_3228_n3085# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X29 AVDD.t120 VB1.t89 a_2712_1638# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X30 AVDD.t119 VB1.t90 a_2002_1638# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X31 AVSS.t202 IREF.t12 a_11544_2488# AVSS.t191 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X32 VB3.t15 VB1.t91 a_3228_4980# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X33 AVSS.t167 AVSS.t165 AVSS.t167 AVSS.t166 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X34 AVDD.t418 AVDD.t417 AVDD.t418 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X35 a_1486_6484# VB1.t92 AVDD.t118 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X36 VB1.t70 VB1.t69 a_3228_2103# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X37 AVSS.t164 AVSS.t163 AVSS.t164 AVSS.t37 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X38 a_11544_2488# IREF.t13 VB1.t1 AVSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X39 a_1486_n77# VB1.t93 AVDD.t117 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X40 a_4970_4093# VB1.t94 VB3.t31 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X41 AVDD.t416 AVDD.t415 AVDD.t416 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X42 AVSS.t162 AVSS.t160 AVSS.t162 AVSS.t161 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X43 AVDD.t116 VB1.t95 a_3744_n2468# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X44 AVDD.t414 AVDD.t412 AVDD.t413 AVDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X45 a_2002_n964# VB1.t96 VB2.t38 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X46 a_3228_n77# VB1.t97 AVDD.t115 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X47 AVSS.t159 AVSS.t156 AVSS.t158 AVSS.t157 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X48 AVSS.t204 IREF.t14 a_11544_1583# AVSS.t191 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X49 VB2.t44 VB1.t98 a_4454_n2468# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X50 a_2002_2724# VB1.t17 VB1.t18 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X51 AVDD.t114 VB1.t99 a_2712_n2468# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X52 a_3228_n3085# VB1.t100 AVDD.t110 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X53 AVDD.t411 AVDD.t410 AVDD.t411 AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X54 AVDD.t409 AVDD.t407 AVDD.t408 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X55 a_3228_5597# VB1.t101 AVDD.t113 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X56 a_1486_n3085# VB1.t102 AVDD.t112 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X57 AVDD.t406 AVDD.t405 AVDD.t406 AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X58 VB2.t36 VB1.t103 a_1486_n964# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X59 AVDD.t404 AVDD.t403 AVDD.t404 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X60 a_2712_3472# VB1.t104 VB3.t29 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X61 a_8985_205# IREF.t15 AVSS.t206 AVSS.t185 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X62 a_11544_1583# IREF.t0 IREF.t1 AVSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X63 a_2712_542# VB1.t67 VB1.t68 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X64 VB1.t60 VB1.t59 a_1486_2724# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X65 AVDD.t402 AVDD.t401 AVDD.t402 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X66 a_3228_1638# VB1.t105 AVDD.t111 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X67 a_8985_2488# VB2.t46 AVSS.t201 AVSS.t185 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X68 AVSS.t155 AVSS.t153 AVSS.t155 AVSS.t154 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X69 a_1486_n964# VB1.t106 AVDD.t109 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X70 AVDD.t400 AVDD.t398 AVDD.t399 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X71 a_2002_n2468# VB1.t107 VB2.t37 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X72 AVSS.t152 AVSS.t149 AVSS.t151 AVSS.t150 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X73 AVDD.t108 VB1.t108 a_3744_n77# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X74 a_1486_2724# VB1.t109 AVDD.t107 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X75 a_4970_542# VB1.t55 VB1.t56 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X76 a_2712_n2468# VB1.t110 VB3.t13 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X77 AVDD.t106 VB1.t111 a_4970_4093# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X78 AVDD.t397 AVDD.t396 AVDD.t397 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X79 AVSS.t148 AVSS.t145 AVSS.t147 AVSS.t146 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X80 AVDD.t395 AVDD.t393 AVDD.t394 AVDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X81 AVDD.t392 AVDD.t391 AVDD.t392 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X82 a_8985_1583# VB2.t47 AVSS.t200 AVSS.t185 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X83 AVDD.t390 AVDD.t388 AVDD.t389 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X84 AVDD.t387 AVDD.t386 AVDD.t387 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X85 AVDD.t385 AVDD.t384 AVDD.t385 AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X86 AVSS.t144 AVSS.t143 AVSS.t144 AVSS.t59 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X87 AVDD.t383 AVDD.t382 AVDD.t383 AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X88 a_4970_3472# VB1.t112 VB2.t6 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X89 AVDD.t381 AVDD.t380 AVDD.t381 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X90 AVDD.t379 AVDD.t378 AVDD.t379 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X91 a_10519_6762# VB4.t17 AVDD.t6 AVDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X92 AVSS.t199 VB2.t48 a_11544_205# AVSS.t191 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X93 AVDD.t377 AVDD.t375 AVDD.t376 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X94 IREF.t7 IREF.t6 a_8985_1111# AVSS.t184 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X95 AVDD.t105 VB1.t113 a_2712_1009# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X96 AVDD.t104 VB1.t114 a_2002_1009# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X97 AVDD.t374 AVDD.t372 AVDD.t373 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X98 AVDD.t371 AVDD.t369 AVDD.t370 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X99 AVDD.t368 AVDD.t366 AVDD.t367 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X100 AVSS.t142 AVSS.t140 AVSS.t141 AVSS.t48 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X101 a_1486_542# VB1.t115 AVDD.t103 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X102 AVDD.t365 AVDD.t363 AVDD.t364 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X103 a_3228_542# VB1.t116 AVDD.t101 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X104 AVDD.t362 AVDD.t360 AVDD.t361 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X105 VB3.t36 VB3.t35 a_10086_n3072# AVSS.t37 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X106 AVSS.t139 AVSS.t137 AVSS.t138 AVSS.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X107 AVSS.t136 AVSS.t134 AVSS.t135 AVSS.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X108 VB2.t33 VB1.t117 a_4454_6484# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X109 a_10691_2488# VB2.t49 AVSS.t198 AVSS.t188 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X110 AVSS.t133 AVSS.t131 AVSS.t133 AVSS.t132 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X111 a_2002_4980# VB1.t118 VB2.t35 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X112 AVSS.t130 AVSS.t128 AVSS.t129 AVSS.t85 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X113 a_4454_6484# VB1.t119 AVDD.t102 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X114 VB4.t7 VB4.t6 a_10777_5228# AVDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X115 AVDD.t359 AVDD.t358 AVDD.t359 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X116 AVDD.t100 VB1.t120 a_4970_3472# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X117 AVDD.t357 AVDD.t355 AVDD.t356 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X118 a_2002_2103# VB1.t63 VB1.t64 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X119 AVDD.t354 AVDD.t352 AVDD.t353 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X120 AVDD.t99 VB1.t121 a_4970_n1581# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X121 VB2.t39 VB1.t122 a_1486_4980# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X122 VB2.t41 VB1.t123 a_3228_n1581# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X123 AVSS.t127 AVSS.t124 AVSS.t126 AVSS.t125 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X124 AVDD.t98 VB1.t124 a_3744_542# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X125 a_3228_1009# VB1.t125 AVDD.t97 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X126 a_10691_1583# VB2.t50 AVSS.t197 AVSS.t188 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X127 AVSS.t187 IREF.t16 a_9838_2488# AVSS.t182 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X128 a_10777_5228# VB4.t18 a_10519_5228# AVDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X129 AVSS.t123 AVSS.t121 AVSS.t122 AVSS.t48 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X130 VB1.t32 VB1.t31 a_1486_2103# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X131 AVDD.t351 AVDD.t349 AVDD.t350 AVDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X132 VB2.t40 VB1.t126 a_4454_n964# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X133 a_1486_4980# VB1.t127 AVDD.t96 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X134 AVDD.t348 AVDD.t346 AVDD.t347 AVDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X135 VB1.t62 VB1.t61 a_4454_2724# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X136 AVDD.t345 AVDD.t344 AVDD.t345 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X137 AVSS.t183 IREF.t17 a_9838_1583# AVSS.t182 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X138 AVDD.t343 AVDD.t342 AVDD.t343 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X139 a_1486_2103# VB1.t128 AVDD.t95 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X140 AVDD.t94 VB1.t129 a_2712_4093# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X141 AVDD.t93 VB1.t130 a_2002_4093# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X142 a_4454_n964# VB1.t131 AVDD.t92 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X143 a_3228_n1581# VB1.t132 AVDD.t91 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X144 a_4454_2724# VB1.t133 AVDD.t90 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X145 AVDD.t341 AVDD.t339 AVDD.t340 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X146 a_1486_n1581# VB1.t134 AVDD.t89 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X147 AVSS.t120 AVSS.t119 AVSS.t120 AVSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X148 AVDD.t338 AVDD.t336 AVDD.t337 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X149 AVDD.t335 AVDD.t334 AVDD.t335 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X150 AVSS.t196 VB2.t51 a_8132_1111# AVSS.t180 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X151 AVDD.t88 VB1.t135 a_3744_5597# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X152 AVSS.t118 AVSS.t117 AVSS.t118 AVSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X153 a_9570_n3072# VB3.t37 AVSS.t6 AVSS.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X154 AVSS.t116 AVSS.t114 AVSS.t115 AVSS.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X155 AVDD.t333 AVDD.t331 AVDD.t332 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X156 AVDD.t330 AVDD.t329 AVDD.t330 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X157 AVDD.t328 AVDD.t326 AVDD.t327 AVDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X158 AVDD.t87 VB1.t136 a_3744_1638# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X159 AVDD.t325 AVDD.t323 AVDD.t324 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X160 a_3744_5597# VB1.t137 VB2.t11 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X161 AVSS.t113 AVSS.t111 AVSS.t112 AVSS.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X162 AVDD.t322 AVDD.t320 AVDD.t321 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X163 a_3228_4093# VB1.t138 AVDD.t86 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X164 AVSS.t110 AVSS.t108 AVSS.t110 AVSS.t109 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X165 a_3744_1638# VB1.t71 VB1.t72 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X166 VB2.t1 VB1.t139 a_3228_5597# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X167 VB1.t3 IREF.t18 a_10691_205# AVSS.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X168 AVDD.t85 VB1.t140 a_2712_3472# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X169 AVDD.t84 VB1.t141 a_2002_3472# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X170 AVDD.t319 AVDD.t317 AVDD.t318 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X171 AVDD.t316 AVDD.t314 AVDD.t315 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X172 AVDD.t313 AVDD.t311 AVDD.t312 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X173 VB1.t58 VB1.t57 a_3228_1638# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X174 a_3744_n3085# VB1.t142 VB2.t8 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X175 a_4454_n3085# VB1.t143 AVDD.t83 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X176 VB2.t43 VB1.t144 a_4454_4980# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X177 a_3744_n77# VB1.t145 VB2.t4 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X178 AVDD.t310 AVDD.t309 AVDD.t310 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X179 VB4.t1 VB4.t0 a_10777_6762# AVDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X180 a_2712_6484# VB1.t146 VB3.t17 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X181 VB1.t12 VB1.t11 a_4454_2103# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X182 a_4454_4980# VB1.t147 AVDD.t82 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X183 AVDD.t308 AVDD.t306 AVDD.t307 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X184 AVDD.t305 AVDD.t303 AVDD.t304 AVDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X185 AVDD.t302 AVDD.t300 AVDD.t301 AVDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X186 a_10777_6762# VB4.t19 a_10519_6762# AVDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X187 a_10519_5531# VB4.t20 AVDD.t5 AVDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X188 a_11544_205# VB2.t52 VB4.t13 AVSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X189 a_4454_2103# VB1.t148 AVDD.t81 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X190 a_3228_3472# VB1.t149 AVDD.t80 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X191 VB3.t25 VB1.t150 a_1486_n3085# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X192 AVDD.t299 AVDD.t298 AVDD.t299 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X193 AVDD.t297 AVDD.t296 AVDD.t297 AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X194 AVSS.t107 AVSS.t105 AVSS.t107 AVSS.t106 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X195 AVDD.t295 AVDD.t293 AVDD.t294 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X196 AVDD.t79 VB1.t151 a_3744_1009# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X197 a_4970_6484# VB1.t152 VB2.t16 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X198 AVSS.t104 AVSS.t103 AVSS.t104 AVSS.t59 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X199 AVDD.t292 AVDD.t291 AVDD.t292 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X200 a_2712_n964# VB1.t153 VB3.t1 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X201 a_2712_2724# VB1.t43 VB1.t44 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X202 AVSS.t102 AVSS.t100 AVSS.t101 AVSS.t85 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X203 VB4.t14 VB2.t53 a_8985_2488# AVSS.t184 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X204 a_3744_1009# VB1.t53 VB1.t54 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X205 AVSS.t99 AVSS.t97 AVSS.t98 AVSS.t48 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X206 AVDD.t290 AVDD.t289 AVDD.t290 AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X207 AVDD.t288 AVDD.t287 AVDD.t288 AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X208 AVSS.t96 AVSS.t95 AVSS.t96 AVSS.t59 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X209 a_3744_542# VB1.t73 VB1.t74 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X210 VB1.t16 VB1.t15 a_3228_1009# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X211 VB2.t25 VB2.t24 a_8985_1583# AVSS.t184 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X212 AVDD.t286 AVDD.t285 AVDD.t286 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X213 AVSS.t94 AVSS.t92 AVSS.t93 AVSS.t48 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X214 AVDD.t284 AVDD.t283 AVDD.t284 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X215 a_2002_5597# VB1.t154 VB3.t2 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X216 a_4970_n964# VB1.t155 VB2.t30 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X217 AVDD.t282 AVDD.t281 AVDD.t282 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X218 AVSS.t91 AVSS.t90 AVSS.t91 AVSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X219 AVDD.t280 AVDD.t278 AVDD.t279 AVDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X220 a_4970_2724# VB1.t41 VB1.t42 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X221 AVDD.t78 VB1.t156 a_4970_6484# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X222 AVDD.t77 VB1.t157 a_4970_n2468# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X223 a_2002_1638# VB1.t7 VB1.t8 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X224 VB3.t23 VB1.t158 a_3228_n2468# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X225 AVSS.t195 VB2.t54 a_9838_205# AVSS.t182 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X226 VB3.t19 VB1.t159 a_1486_5597# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X227 a_8132_205# VB2.t55 VB4.t11 AVSS.t194 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X228 AVDD.t277 AVDD.t276 AVDD.t277 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X229 VB1.t26 VB1.t25 a_1486_1638# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X230 AVDD.t12 VB1.t160 a_3744_4093# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X231 a_1486_5597# VB1.t161 AVDD.t76 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X232 AVDD.t275 AVDD.t274 AVDD.t275 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X233 AVSS.t89 AVSS.t88 AVSS.t89 AVSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X234 AVDD.t273 AVDD.t272 AVDD.t273 AVDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X235 AVDD.t271 AVDD.t270 AVDD.t271 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X236 AVDD.t269 AVDD.t268 AVDD.t269 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X237 a_3744_n1581# VB1.t162 VB2.t5 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X238 a_10691_205# IREF.t19 AVSS.t203 AVSS.t188 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X239 AVDD.t267 AVDD.t265 AVDD.t266 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X240 AVDD.t74 VB1.t163 a_2712_n77# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X241 a_1486_1638# VB1.t164 AVDD.t75 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X242 AVDD.t73 VB1.t165 a_4970_n964# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X243 a_4454_n1581# VB1.t166 AVDD.t72 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X244 a_3228_n2468# VB1.t167 AVDD.t71 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X245 VB3.t22 VB1.t168 a_4454_n77# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X246 a_3744_4093# VB1.t169 VB2.t13 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X247 AVDD.t264 AVDD.t263 AVDD.t264 AVDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X248 a_1486_n2468# VB1.t170 AVDD.t70 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X249 AVSS.t87 AVSS.t84 AVSS.t86 AVSS.t85 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X250 AVDD.t69 VB1.t171 a_4970_2724# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X251 AVDD.t68 VB1.t172 a_2002_n3085# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X252 a_2712_4980# VB1.t173 VB3.t28 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X253 AVSS.t83 AVSS.t81 AVSS.t83 AVSS.t82 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X254 VB2.t2 VB1.t174 a_3228_4093# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X255 AVSS.t205 IREF.t20 a_8132_2488# AVSS.t180 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X256 a_2712_2103# VB1.t39 VB1.t40 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X257 VB3.t11 VB1.t175 a_1486_n1581# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X258 AVDD.t262 AVDD.t260 AVDD.t261 AVDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X259 AVDD.t259 AVDD.t257 AVDD.t258 AVDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X260 AVDD.t256 AVDD.t255 AVDD.t256 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X261 AVSS.t181 IREF.t21 a_8132_1583# AVSS.t180 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X262 AVDD.t67 VB1.t176 a_3744_3472# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X263 AVDD.t254 AVDD.t253 AVDD.t254 AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X264 a_4970_4980# VB1.t177 VB2.t15 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X265 VB2.t32 VB1.t178 a_3228_n77# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X266 a_2002_1009# VB1.t49 VB1.t50 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X267 AVDD.t66 VB1.t179 a_4970_n77# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X268 AVDD.t65 VB1.t180 a_2002_6484# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X269 AVDD.t64 VB1.t181 a_2712_6484# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X270 a_4970_2103# VB1.t9 VB1.t10 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X271 AVDD.t252 AVDD.t251 AVDD.t252 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X272 VB4.t5 VB4.t4 a_10777_5531# AVDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X273 AVDD.t250 AVDD.t249 AVDD.t250 AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X274 a_3744_3472# VB1.t182 VB3.t21 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X275 AVDD.t248 AVDD.t246 AVDD.t247 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X276 a_4970_n3085# VB1.t183 VB3.t6 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X277 a_2002_n77# VB1.t184 VB3.t14 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X278 VB1.t38 VB1.t37 a_1486_1009# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X279 AVDD.t63 VB1.t185 a_2712_542# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X280 AVDD.t245 AVDD.t243 AVDD.t244 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X281 a_10777_5531# VB4.t21 a_10519_5531# AVDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X282 VB1.t34 VB1.t33 a_4454_542# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X283 AVDD.t242 AVDD.t240 AVDD.t241 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X284 AVDD.t239 AVDD.t237 AVDD.t238 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X285 VB1.t2 IREF.t22 a_8985_205# AVSS.t184 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X286 VB3.t7 VB1.t186 a_3228_3472# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X287 VB3.t33 VB1.t187 a_4454_5597# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X288 AVDD.t236 AVDD.t235 AVDD.t236 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X289 AVDD.t234 AVDD.t233 AVDD.t234 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X290 a_1486_1009# VB1.t188 AVDD.t62 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X291 AVDD.t232 AVDD.t231 AVDD.t232 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X292 VB1.t36 VB1.t35 a_4454_1638# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X293 AVDD.t230 AVDD.t229 AVDD.t230 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X294 a_4454_5597# VB1.t189 AVDD.t61 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X295 AVDD.t60 VB1.t190 a_3744_n3085# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X296 AVDD.t59 VB1.t191 a_4970_4980# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X297 IREF.t3 IREF.t2 a_10691_1111# AVSS.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X298 AVDD.t228 AVDD.t226 AVDD.t227 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X299 AVDD.t58 VB1.t192 a_2712_n964# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X300 AVDD.t57 VB1.t193 a_2002_n964# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X301 AVDD.t225 AVDD.t223 AVDD.t224 AVDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X302 VB3.t10 VB1.t194 a_4454_n3085# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X303 AVDD.t56 VB1.t195 a_2712_2724# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X304 AVDD.t55 VB1.t196 a_2002_2724# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X305 a_3228_6484# VB1.t197 AVDD.t54 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X306 AVDD.t53 VB1.t198 a_2712_n3085# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X307 AVDD.t222 AVDD.t221 AVDD.t222 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X308 a_4454_1638# VB1.t199 AVDD.t52 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X309 AVDD.t51 VB1.t200 a_4970_2103# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X310 AVDD.t220 AVDD.t218 AVDD.t219 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X311 AVSS.t80 AVSS.t79 AVSS.t80 AVSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X312 AVSS.t78 AVSS.t76 AVSS.t77 AVSS.t33 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X313 a_10519_5995# VB4.t22 AVDD.t4 AVDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X314 AVSS.t75 AVSS.t73 AVSS.t74 AVSS.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X315 VB1.t46 VB1.t45 a_3228_542# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X316 AVDD.t50 VB1.t201 a_4970_542# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X317 a_2002_4093# VB1.t202 VB3.t12 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X318 a_2002_n3085# VB1.t203 VB3.t3 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X319 AVDD.t217 AVDD.t216 AVDD.t217 AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X320 AVSS.t72 AVSS.t71 AVSS.t72 AVSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X321 AVSS.t70 AVSS.t68 AVSS.t70 AVSS.t69 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X322 AVDD.t215 AVDD.t213 AVDD.t214 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X323 a_2712_n3085# VB1.t204 VB2.t14 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X324 AVDD.t212 AVDD.t211 AVDD.t212 AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X325 AVDD.t210 AVDD.t209 AVDD.t210 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X326 AVDD.t208 AVDD.t207 AVDD.t208 AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X327 AVDD.t10 VB1.t205 a_2002_n1581# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X328 a_2002_542# VB1.t27 VB1.t28 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X329 VB3.t32 VB1.t206 a_1486_4093# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X330 a_3228_n964# VB1.t207 AVDD.t49 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X331 a_8132_1111# VB2.t26 VB2.t27 AVSS.t194 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X332 a_3228_2724# VB1.t208 AVDD.t48 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X333 AVDD.t206 AVDD.t204 AVDD.t205 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X334 AVDD.t203 AVDD.t201 AVDD.t202 AVDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X335 a_9838_1111# VB2.t20 VB2.t21 AVSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X336 a_1486_4093# VB1.t209 AVDD.t47 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X337 AVDD.t200 AVDD.t199 AVDD.t200 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X338 AVSS.t67 AVSS.t66 AVSS.t67 AVSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X339 AVDD.t198 AVDD.t197 AVDD.t198 AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X340 AVDD.t196 AVDD.t195 AVDD.t196 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X341 AVDD.t194 AVDD.t191 AVDD.t193 AVDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X342 AVDD.t190 AVDD.t188 AVDD.t189 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X343 AVDD.t187 AVDD.t185 AVDD.t186 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X344 VB1.t22 VB1.t21 a_4454_1009# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X345 AVSS.t193 VB2.t56 a_8132_205# AVSS.t180 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X346 AVDD.t184 AVDD.t182 AVDD.t183 AVDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X347 AVSS.t65 AVSS.t64 AVSS.t65 AVSS.t59 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X348 a_4454_n77# VB1.t210 AVDD.t46 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X349 AVDD.t181 AVDD.t180 AVDD.t181 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X350 AVDD.t179 AVDD.t177 AVDD.t178 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X351 a_2002_3472# VB1.t211 VB2.t29 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X352 AVSS.t63 AVSS.t61 AVSS.t63 AVSS.t62 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X353 AVDD.t45 VB1.t212 a_2712_4980# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X354 AVDD.t44 VB1.t213 a_2002_4980# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X355 a_4454_1009# VB1.t214 AVDD.t43 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X356 AVSS.t60 AVSS.t58 AVSS.t60 AVSS.t59 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X357 AVDD.t176 AVDD.t174 AVDD.t175 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X358 AVSS.t57 AVSS.t55 AVSS.t56 AVSS.t48 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X359 AVDD.t173 AVDD.t172 AVDD.t173 AVDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X360 a_4970_n1581# VB1.t215 VB3.t16 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X361 a_3744_n2468# VB1.t216 VB3.t30 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X362 AVDD.t42 VB1.t217 a_2712_2103# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X363 AVDD.t41 VB1.t218 a_2002_2103# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X364 VB2.t12 VB1.t219 a_1486_3472# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X365 AVSS.t192 VB2.t57 a_11544_1111# AVSS.t191 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X366 a_4454_n2468# VB1.t220 AVDD.t40 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X367 AVSS.t54 AVSS.t51 AVSS.t53 AVSS.t52 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X368 AVSS.t50 AVSS.t47 AVSS.t49 AVSS.t48 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X369 AVDD.t171 AVDD.t170 AVDD.t171 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X370 a_10086_n3072# VB3.t38 a_9828_n3072# AVSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X371 AVDD.t169 AVDD.t168 AVDD.t169 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X372 AVDD.t167 AVDD.t166 AVDD.t167 AVDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X373 a_1486_3472# VB1.t221 AVDD.t39 AVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X374 a_2712_5597# VB1.t222 VB2.t3 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X375 AVDD.t165 AVDD.t164 AVDD.t165 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X376 a_11544_1111# VB2.t22 VB2.t23 AVSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X377 a_10519_6298# VB4.t23 AVDD.t3 AVDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X378 AVDD.t37 VB1.t223 a_3744_n1581# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X379 AVDD.t163 AVDD.t161 AVDD.t162 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X380 AVDD.t160 AVDD.t158 AVDD.t159 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X381 a_2712_1638# VB1.t19 VB1.t20 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X382 VB3.t34 VB1.t224 a_4454_n1581# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X383 AVDD.t157 AVDD.t155 AVDD.t156 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X384 AVDD.t36 VB1.t225 a_2712_n1581# AVDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X385 VB2.t17 VB1.t226 a_1486_n2468# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X386 a_3228_4980# VB1.t227 AVDD.t34 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X387 AVSS.t46 AVSS.t43 AVSS.t45 AVSS.t44 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X388 a_9828_n3072# VB3.t39 a_9570_n3072# AVSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X389 a_3228_2103# VB1.t228 AVDD.t33 AVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X390 a_8985_1111# IREF.t23 AVSS.t186 AVSS.t185 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X391 VB3.t5 VB1.t229 a_1486_n77# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X392 VB3.t9 VB1.t230 a_4454_4093# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X393 AVDD.t31 VB1.t231 a_3744_6484# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X394 AVSS.t42 AVSS.t39 AVSS.t41 AVSS.t40 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X395 AVSS.t38 AVSS.t36 AVSS.t38 AVSS.t37 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X396 a_4454_542# VB1.t232 AVDD.t30 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X397 a_4970_5597# VB1.t233 VB3.t8 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X398 a_2002_n1581# VB1.t234 VB3.t0 AVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X399 a_4454_4093# VB1.t235 AVDD.t28 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X400 AVDD.t154 AVDD.t152 AVDD.t153 AVDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X401 a_3744_6484# VB1.t236 VB3.t24 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X402 a_2712_n1581# VB1.t237 VB2.t42 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X403 a_4970_1638# VB1.t29 VB1.t30 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X404 AVDD.t26 VB1.t238 a_2002_n77# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X405 VB4.t3 VB4.t2 a_10777_5995# AVDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X406 VB3.t26 VB1.t239 a_3228_6484# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X407 AVSS.t35 AVSS.t32 AVSS.t34 AVSS.t33 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X408 AVDD.t151 AVDD.t148 AVDD.t150 AVDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X409 AVDD.t13 VB1.t240 a_3744_n964# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X410 a_10777_5995# VB4.t24 a_10519_5995# AVDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X411 AVDD.t147 AVDD.t146 AVDD.t147 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X412 AVDD.t25 VB1.t241 a_3744_2724# AVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X413 AVDD.t145 AVDD.t143 AVDD.t145 AVDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X414 AVSS.t31 AVSS.t29 AVSS.t31 AVSS.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X415 AVDD.t24 VB1.t242 a_4970_5597# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X416 AVDD.t142 AVDD.t140 AVDD.t142 AVDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X417 VB4.t12 VB2.t58 a_10691_2488# AVSS.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X418 AVDD.t139 AVDD.t137 AVDD.t138 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X419 a_3744_n964# VB1.t243 VB3.t20 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X420 VB2.t10 VB1.t244 a_4454_3472# AVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X421 AVDD.t136 AVDD.t133 AVDD.t135 AVDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X422 a_3744_2724# VB1.t23 VB1.t24 AVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X423 a_10691_1111# IREF.t24 AVSS.t189 AVSS.t188 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X424 AVSS.t28 AVSS.t25 AVSS.t27 AVSS.t26 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X425 AVDD.t21 VB1.t245 a_4970_1638# AVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X426 AVSS.t24 AVSS.t23 AVSS.t24 AVSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X427 a_2712_1009# VB1.t51 VB1.t52 AVDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X428 VB1.t48 VB1.t47 a_1486_542# AVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X429 VB3.t18 VB1.t246 a_3228_n964# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X430 a_4454_3472# VB1.t247 AVDD.t17 AVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X431 VB2.t19 VB2.t18 a_10691_1583# AVSS.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X432 VB1.t14 VB1.t13 a_3228_2724# AVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X433 AVSS.t22 AVSS.t21 AVSS.t22 AVSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X434 AVSS.t20 AVSS.t17 AVSS.t19 AVSS.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X435 AVSS.t190 VB2.t59 a_9838_1111# AVSS.t182 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X436 AVDD.t132 AVDD.t129 AVDD.t131 AVDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X437 AVSS.t16 AVSS.t14 AVSS.t16 AVSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X438 AVSS.t13 AVSS.t11 AVSS.t12 AVSS.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X439 AVSS.t10 AVSS.t7 AVSS.t9 AVSS.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X440 AVDD.t14 VB1.t248 a_2002_542# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X441 AVDD.t128 AVDD.t127 AVDD.t128 AVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X442 AVDD.t9 VB1.t249 a_2002_n2468# AVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
R0 VB2.n45 VB2.t3 235.565
R1 VB2.n52 VB2.t0 235.565
R2 VB2.n59 VB2.t9 235.565
R3 VB2.n68 VB2.t42 235.565
R4 VB2.n62 VB2.t14 235.565
R5 VB2.n65 VB2.n63 210.161
R6 VB2.n43 VB2.n41 210.157
R7 VB2.n49 VB2.n47 210.157
R8 VB2.n56 VB2.n54 210.157
R9 VB2.n73 VB2.n71 210.15
R10 VB2.n45 VB2.n44 205.238
R11 VB2.n52 VB2.n51 205.238
R12 VB2.n59 VB2.n58 205.238
R13 VB2.n68 VB2.n67 205.238
R14 VB2.n62 VB2.n61 205.238
R15 VB2.n73 VB2.n72 204.861
R16 VB2.n65 VB2.n64 204.859
R17 VB2.n43 VB2.n42 204.857
R18 VB2.n49 VB2.n48 204.857
R19 VB2.n56 VB2.n55 204.857
R20 VB2.n17 VB2.t47 114.496
R21 VB2.n81 VB2.t55 114.496
R22 VB2.n101 VB2.t48 114.496
R23 VB2.n9 VB2.t46 114.468
R24 VB2.n110 VB2.t57 114.466
R25 VB2.n2 VB2.t58 114.466
R26 VB2.n11 VB2.t53 103.459
R27 VB2.n4 VB2.t49 103.459
R28 VB2.n19 VB2.t24 103.459
R29 VB2.n36 VB2.t50 103.459
R30 VB2.n28 VB2.t18 103.459
R31 VB2.n138 VB2.t20 103.459
R32 VB2.n146 VB2.t59 103.459
R33 VB2.n124 VB2.t26 103.459
R34 VB2.n132 VB2.t51 103.459
R35 VB2.n112 VB2.t22 103.459
R36 VB2.n83 VB2.t56 103.459
R37 VB2.n88 VB2.t45 103.459
R38 VB2.n96 VB2.t54 103.459
R39 VB2.n103 VB2.t52 103.459
R40 VB2.n21 VB2.t25 87.5271
R41 VB2.n26 VB2.t19 87.5245
R42 VB2.n122 VB2.t27 87.4861
R43 VB2.n137 VB2.t21 87.4848
R44 VB2.n114 VB2.t23 87.4826
R45 VB2.n41 VB2.t31 28.5655
R46 VB2.n41 VB2.t28 28.5655
R47 VB2.n42 VB2.t16 28.5655
R48 VB2.n42 VB2.t33 28.5655
R49 VB2.n44 VB2.t11 28.5655
R50 VB2.n44 VB2.t1 28.5655
R51 VB2.n47 VB2.t35 28.5655
R52 VB2.n47 VB2.t39 28.5655
R53 VB2.n48 VB2.t15 28.5655
R54 VB2.n48 VB2.t43 28.5655
R55 VB2.n51 VB2.t13 28.5655
R56 VB2.n51 VB2.t2 28.5655
R57 VB2.n54 VB2.t29 28.5655
R58 VB2.n54 VB2.t12 28.5655
R59 VB2.n55 VB2.t6 28.5655
R60 VB2.n55 VB2.t10 28.5655
R61 VB2.n58 VB2.t4 28.5655
R62 VB2.n58 VB2.t32 28.5655
R63 VB2.n67 VB2.t5 28.5655
R64 VB2.n67 VB2.t41 28.5655
R65 VB2.n63 VB2.t37 28.5655
R66 VB2.n63 VB2.t17 28.5655
R67 VB2.n64 VB2.t7 28.5655
R68 VB2.n64 VB2.t44 28.5655
R69 VB2.n61 VB2.t8 28.5655
R70 VB2.n61 VB2.t34 28.5655
R71 VB2.n72 VB2.t30 28.5655
R72 VB2.n72 VB2.t40 28.5655
R73 VB2.n71 VB2.t38 28.5655
R74 VB2.n71 VB2.t36 28.5655
R75 VB2.n12 VB2.n11 21.9607
R76 VB2.n11 VB2.n10 21.9607
R77 VB2.n4 VB2.n3 21.9607
R78 VB2.n5 VB2.n4 21.9607
R79 VB2.n20 VB2.n19 21.9607
R80 VB2.n19 VB2.n18 21.9607
R81 VB2.n36 VB2.n35 21.9607
R82 VB2.n37 VB2.n36 21.9607
R83 VB2.n28 VB2.n27 21.9607
R84 VB2.n29 VB2.n28 21.9607
R85 VB2.n138 VB2.n136 21.9607
R86 VB2.n139 VB2.n138 21.9607
R87 VB2.n147 VB2.n146 21.9607
R88 VB2.n146 VB2.n145 21.9607
R89 VB2.n124 VB2.n123 21.9607
R90 VB2.n125 VB2.n124 21.9607
R91 VB2.n133 VB2.n132 21.9607
R92 VB2.n132 VB2.n131 21.9607
R93 VB2.n112 VB2.n111 21.9607
R94 VB2.n113 VB2.n112 21.9607
R95 VB2.n84 VB2.n83 21.9607
R96 VB2.n83 VB2.n82 21.9607
R97 VB2.n88 VB2.n87 21.9607
R98 VB2.n89 VB2.n88 21.9607
R99 VB2.n97 VB2.n96 21.9607
R100 VB2.n96 VB2.n95 21.9607
R101 VB2.n103 VB2.n102 21.9607
R102 VB2.n104 VB2.n103 21.9607
R103 VB2.n75 VB2.n74 5.80879
R104 VB2.n31 VB2.n26 4.61479
R105 VB2.n127 VB2.n122 4.61479
R106 VB2.n85 VB2.n84 4.51108
R107 VB2.n89 VB2.n86 4.51108
R108 VB2.n105 VB2.n104 4.51012
R109 VB2.n98 VB2.n97 4.50819
R110 VB2.n38 VB2.n37 4.50723
R111 VB2.n13 VB2.n12 4.50541
R112 VB2.n134 VB2.n133 4.50539
R113 VB2.n148 VB2.n147 4.50406
R114 VB2.n6 VB2.n5 4.50363
R115 VB2.n8 VB2.n7 4.5005
R116 VB2.n1 VB2.n0 4.5005
R117 VB2.n16 VB2.n15 4.5005
R118 VB2.n22 VB2.n21 4.5005
R119 VB2.n24 VB2.n23 4.5005
R120 VB2.n34 VB2.n33 4.5005
R121 VB2.n32 VB2.n25 4.5005
R122 VB2.n31 VB2.n30 4.5005
R123 VB2.n127 VB2.n126 4.5005
R124 VB2.n128 VB2.n121 4.5005
R125 VB2.n130 VB2.n129 4.5005
R126 VB2.n120 VB2.n119 4.5005
R127 VB2.n137 VB2.n135 4.5005
R128 VB2.n141 VB2.n140 4.5005
R129 VB2.n142 VB2.n118 4.5005
R130 VB2.n144 VB2.n143 4.5005
R131 VB2.n117 VB2.n116 4.5005
R132 VB2.n115 VB2.n114 4.5005
R133 VB2.n109 VB2.n108 4.5005
R134 VB2.n91 VB2.n90 4.5005
R135 VB2.n92 VB2.n78 4.5005
R136 VB2.n94 VB2.n93 4.5005
R137 VB2.n77 VB2.n76 4.5005
R138 VB2.n80 VB2.n79 4.5005
R139 VB2.n100 VB2.n99 4.5005
R140 VB2.n66 VB2.n62 4.46199
R141 VB2.n46 VB2.n45 4.29389
R142 VB2.n53 VB2.n52 4.29389
R143 VB2.n60 VB2.n59 4.29389
R144 VB2.n69 VB2.n68 4.29389
R145 VB2.n135 VB2.n134 2.41836
R146 VB2.n86 VB2.n85 2.41836
R147 VB2.n46 VB2.n43 2.17117
R148 VB2.n50 VB2.n49 2.10286
R149 VB2.n57 VB2.n56 2.10286
R150 VB2.n66 VB2.n65 2.10286
R151 VB2.n149 VB2.n115 1.89775
R152 VB2.n106 VB2.n105 1.89739
R153 VB2.n39 VB2.n22 1.88203
R154 VB2.n14 VB2.n13 1.88167
R155 VB2.n2 VB2.n0 1.34982
R156 VB2.n110 VB2.n108 1.34941
R157 VB2.n9 VB2.n7 1.3492
R158 VB2.n101 VB2.n99 1.33272
R159 VB2.n17 VB2.n15 1.33239
R160 VB2.n81 VB2.n79 1.33239
R161 VB2.n40 VB2.n14 1.13717
R162 VB2.n74 VB2.n70 1.09471
R163 VB2.n107 VB2.n106 1.09471
R164 VB2.n150 VB2.n149 1.09471
R165 VB2.n40 VB2.n39 1.09471
R166 VB2.n74 VB2.n73 0.996725
R167 VB2.n60 VB2.n57 0.579697
R168 VB2.n14 VB2.n6 0.379888
R169 VB2.n39 VB2.n38 0.379529
R170 VB2.n106 VB2.n98 0.364174
R171 VB2.n149 VB2.n148 0.363815
R172 VB2.n75 VB2 0.225787
R173 VB2.n107 VB2.n75 0.198057
R174 VB2.n57 VB2.n53 0.168447
R175 VB2.n50 VB2.n46 0.16782
R176 VB2.n33 VB2.n32 0.166571
R177 VB2.n143 VB2.n142 0.166571
R178 VB2.n129 VB2.n128 0.166571
R179 VB2.n93 VB2.n92 0.166571
R180 VB2.n70 VB2.n69 0.16594
R181 VB2.n102 VB2.n101 0.139606
R182 VB2.n18 VB2.n17 0.138972
R183 VB2.n82 VB2.n81 0.138972
R184 VB2.n13 VB2.n7 0.114786
R185 VB2.n6 VB2.n0 0.114786
R186 VB2.n22 VB2.n15 0.114786
R187 VB2.n32 VB2.n31 0.114786
R188 VB2.n33 VB2.n23 0.114786
R189 VB2.n38 VB2.n23 0.114786
R190 VB2.n148 VB2.n116 0.114786
R191 VB2.n143 VB2.n116 0.114786
R192 VB2.n142 VB2.n141 0.114786
R193 VB2.n141 VB2.n135 0.114786
R194 VB2.n134 VB2.n119 0.114786
R195 VB2.n129 VB2.n119 0.114786
R196 VB2.n128 VB2.n127 0.114786
R197 VB2.n115 VB2.n108 0.114786
R198 VB2.n98 VB2.n76 0.114786
R199 VB2.n93 VB2.n76 0.114786
R200 VB2.n92 VB2.n91 0.114786
R201 VB2.n91 VB2.n86 0.114786
R202 VB2.n85 VB2.n79 0.114786
R203 VB2.n105 VB2.n99 0.114786
R204 VB2 VB2.n150 0.0908967
R205 VB2.n34 VB2.n25 0.0899231
R206 VB2.n94 VB2.n78 0.0899231
R207 VB2 VB2.n40 0.0835333
R208 VB2.n69 VB2.n66 0.0706867
R209 VB2.n53 VB2.n50 0.0688067
R210 VB2.n3 VB2.n2 0.067158
R211 VB2.n111 VB2.n110 0.0660552
R212 VB2.n10 VB2.n9 0.0659917
R213 VB2 VB2.n60 0.0575267
R214 VB2.n37 VB2.n24 0.0553077
R215 VB2.n97 VB2.n77 0.0543462
R216 VB2.n104 VB2.n100 0.0524231
R217 VB2.n20 VB2.n16 0.0514615
R218 VB2.n84 VB2.n80 0.0514615
R219 VB2.n90 VB2.n89 0.0514615
R220 VB2.n30 VB2.n27 0.0505
R221 VB2.n35 VB2.n34 0.0476154
R222 VB2.n95 VB2.n94 0.0466538
R223 VB2.n87 VB2.n78 0.0437692
R224 VB2.n150 VB2.n107 0.0429567
R225 VB2.n29 VB2.n25 0.0428077
R226 VB2.n144 VB2.n118 0.0418701
R227 VB2.n130 VB2.n121 0.0418701
R228 VB2.n5 VB2.n1 0.0259464
R229 VB2.n147 VB2.n117 0.025411
R230 VB2.n126 VB2.n125 0.025411
R231 VB2.n113 VB2.n109 0.0245214
R232 VB2.n12 VB2.n8 0.0241607
R233 VB2.n140 VB2.n139 0.0240765
R234 VB2.n133 VB2.n120 0.0240765
R235 VB2.n145 VB2.n144 0.0218523
R236 VB2.n123 VB2.n121 0.0218523
R237 VB2.n136 VB2.n118 0.0205178
R238 VB2.n131 VB2.n130 0.0205178
R239 VB2.n30 VB2.n29 0.0197308
R240 VB2.n18 VB2.n16 0.0187692
R241 VB2.n82 VB2.n80 0.0187692
R242 VB2.n90 VB2.n87 0.0187692
R243 VB2.n102 VB2.n100 0.0178077
R244 VB2.n95 VB2.n77 0.0158846
R245 VB2.n35 VB2.n24 0.0149231
R246 VB2.n70 VB2 0.0124067
R247 VB2.n27 VB2.n26 0.0120385
R248 VB2.n21 VB2.n20 0.0110769
R249 VB2.n10 VB2.n8 0.00898214
R250 VB2.n140 VB2.n136 0.00895196
R251 VB2.n131 VB2.n120 0.00895196
R252 VB2.n111 VB2.n109 0.00850712
R253 VB2.n145 VB2.n117 0.00761744
R254 VB2.n126 VB2.n123 0.00761744
R255 VB2.n3 VB2.n1 0.00719643
R256 VB2.n139 VB2.n137 0.00539324
R257 VB2.n114 VB2.n113 0.0049484
R258 VB2.n125 VB2.n122 0.00405872
R259 VB4.n4 VB4.t1 231.773
R260 VB4.n60 VB4.t5 231.625
R261 VB4.n61 VB4.t7 231.625
R262 VB4.n3 VB4.t9 231.625
R263 VB4.n1 VB4.t3 231.625
R264 VB4.n64 VB4.t15 113.684
R265 VB4.n66 VB4.t18 102.6
R266 VB4.n74 VB4.t6 102.6
R267 VB4.n13 VB4.t17 102.6
R268 VB4.n19 VB4.t19 102.6
R269 VB4.n27 VB4.t0 102.6
R270 VB4.n12 VB4.t23 102.6
R271 VB4.n10 VB4.t16 102.6
R272 VB4.n5 VB4.t8 102.6
R273 VB4.n42 VB4.t22 102.6
R274 VB4.n48 VB4.t24 102.6
R275 VB4.n56 VB4.t2 102.6
R276 VB4.n41 VB4.t20 102.6
R277 VB4.n39 VB4.t21 102.6
R278 VB4.n33 VB4.t4 102.6
R279 VB4.n79 VB4.t14 92.3532
R280 VB4.n81 VB4.t11 91.9848
R281 VB4.n79 VB4.t12 89.3182
R282 VB4.n82 VB4.t13 89.1212
R283 VB4.n81 VB4.t10 88.9381
R284 VB4.n66 VB4.n65 21.9522
R285 VB4.n67 VB4.n66 21.9522
R286 VB4.n75 VB4.n74 21.9522
R287 VB4.n74 VB4.n73 21.9522
R288 VB4.n13 VB4.n11 21.9522
R289 VB4.n14 VB4.n13 21.9522
R290 VB4.n19 VB4.n9 21.9522
R291 VB4.n20 VB4.n19 21.9522
R292 VB4.n28 VB4.n27 21.9522
R293 VB4.n27 VB4.n26 21.9522
R294 VB4.n12 VB4.n11 21.9522
R295 VB4.n14 VB4.n12 21.9522
R296 VB4.n10 VB4.n9 21.9522
R297 VB4.n20 VB4.n10 21.9522
R298 VB4.n28 VB4.n5 21.9522
R299 VB4.n26 VB4.n5 21.9522
R300 VB4.n42 VB4.n40 21.9522
R301 VB4.n43 VB4.n42 21.9522
R302 VB4.n48 VB4.n38 21.9522
R303 VB4.n49 VB4.n48 21.9522
R304 VB4.n57 VB4.n56 21.9522
R305 VB4.n56 VB4.n55 21.9522
R306 VB4.n41 VB4.n40 21.9522
R307 VB4.n43 VB4.n41 21.9522
R308 VB4.n39 VB4.n38 21.9522
R309 VB4.n49 VB4.n39 21.9522
R310 VB4.n57 VB4.n33 21.9522
R311 VB4.n55 VB4.n33 21.9522
R312 VB4.n77 VB4.n76 4.5005
R313 VB4.n62 VB4.n0 4.5005
R314 VB4.n72 VB4.n71 4.5005
R315 VB4.n70 VB4.n63 4.5005
R316 VB4.n69 VB4.n68 4.5005
R317 VB4.n82 VB4.n81 2.71364
R318 VB4.n30 VB4.n29 2.2505
R319 VB4.n6 VB4.n2 2.2505
R320 VB4.n25 VB4.n24 2.2505
R321 VB4.n23 VB4.n7 2.2505
R322 VB4.n22 VB4.n21 2.2505
R323 VB4.n18 VB4.n8 2.2505
R324 VB4.n17 VB4.n16 2.2505
R325 VB4.n58 VB4.n32 2.2505
R326 VB4.n46 VB4.n45 2.2505
R327 VB4.n47 VB4.n37 2.2505
R328 VB4.n51 VB4.n50 2.2505
R329 VB4.n52 VB4.n35 2.2505
R330 VB4.n54 VB4.n53 2.2505
R331 VB4.n36 VB4.n34 2.2505
R332 VB4.n31 VB4.n30 1.40428
R333 VB4.n80 VB4.n79 1.379
R334 VB4.n78 VB4.n77 1.33978
R335 VB4 VB4.n82 1.29212
R336 VB4.n32 VB4.n31 1.28412
R337 VB4.n69 VB4.n64 1.23766
R338 VB4.n45 VB4.n44 1.18823
R339 VB4.n16 VB4.n15 1.18805
R340 VB4.n3 VB4.n1 0.317001
R341 VB4.n61 VB4.n60 0.317001
R342 VB4.n76 VB4.n61 0.293199
R343 VB4.n67 VB4.n64 0.243881
R344 VB4 VB4.n80 0.241767
R345 VB4 VB4.n78 0.226413
R346 VB4.n72 VB4.n63 0.2005
R347 VB4.n4 VB4.n3 0.147813
R348 VB4.n60 VB4.n59 0.147813
R349 VB4.n59 VB4.n1 0.147812
R350 VB4.n71 VB4.n70 0.139114
R351 VB4.n80 VB4 0.1227
R352 VB4.n31 VB4 0.106563
R353 VB4.n24 VB4.n23 0.1005
R354 VB4.n53 VB4.n52 0.1005
R355 VB4.n75 VB4.n62 0.0987143
R356 VB4.n16 VB4.n8 0.0951429
R357 VB4.n45 VB4.n37 0.0951429
R358 VB4.n73 VB4.n72 0.0844286
R359 VB4.n29 VB4.n4 0.0836044
R360 VB4.n59 VB4.n58 0.0836044
R361 VB4.n77 VB4.n0 0.0797079
R362 VB4.n71 VB4.n0 0.0797079
R363 VB4.n70 VB4.n69 0.0797079
R364 VB4.n25 VB4.n7 0.0774231
R365 VB4.n54 VB4.n35 0.0774231
R366 VB4.n18 VB4.n17 0.0733022
R367 VB4.n47 VB4.n46 0.0733022
R368 VB4.n68 VB4.n65 0.0665714
R369 VB4.n68 VB4.n67 0.063
R370 VB4.n30 VB4.n2 0.0576429
R371 VB4.n24 VB4.n2 0.0576429
R372 VB4.n23 VB4.n22 0.0576429
R373 VB4.n22 VB4.n8 0.0576429
R374 VB4.n36 VB4.n32 0.0576429
R375 VB4.n53 VB4.n36 0.0576429
R376 VB4.n52 VB4.n51 0.0576429
R377 VB4.n51 VB4.n37 0.0576429
R378 VB4.n65 VB4.n63 0.0487143
R379 VB4.n28 VB4.n6 0.0382747
R380 VB4.n57 VB4.n34 0.0382747
R381 VB4.n17 VB4.n11 0.0355275
R382 VB4.n46 VB4.n40 0.0355275
R383 VB4.n26 VB4.n25 0.0327802
R384 VB4.n55 VB4.n54 0.0327802
R385 VB4.n73 VB4.n62 0.0308571
R386 VB4.n44 VB4.n40 0.0301133
R387 VB4.n15 VB4.n11 0.0297444
R388 VB4.n21 VB4.n9 0.0259121
R389 VB4.n50 VB4.n38 0.0259121
R390 VB4.n21 VB4.n20 0.0245385
R391 VB4.n50 VB4.n49 0.0245385
R392 VB4.n44 VB4.n43 0.021976
R393 VB4.n15 VB4.n14 0.0213493
R394 VB4.n20 VB4.n18 0.0204176
R395 VB4.n49 VB4.n47 0.0204176
R396 VB4.n9 VB4.n7 0.019044
R397 VB4.n38 VB4.n35 0.019044
R398 VB4.n76 VB4.n75 0.0165714
R399 VB4.n26 VB4.n6 0.0121758
R400 VB4.n55 VB4.n34 0.0121758
R401 VB4.n78 VB4 0.00817667
R402 VB4.n29 VB4.n28 0.00668132
R403 VB4.n58 VB4.n57 0.00668132
R404 AVSS.n516 AVSS.n390 4200.73
R405 AVSS.n647 AVSS.n393 2155.41
R406 AVSS.n1679 AVSS.n1311 2120.65
R407 AVSS.n1682 AVSS.n1681 2045.32
R408 AVSS.n1751 AVSS.n42 2045.32
R409 AVSS.n906 AVSS.n280 1842.53
R410 AVSS.n1754 AVSS.n14 1761.41
R411 AVSS.n873 AVSS.n793 1558.62
R412 AVSS.n1682 AVSS.n1302 585
R413 AVSS.n1685 AVSS.n1684 585
R414 AVSS.n1394 AVSS.n1305 585
R415 AVSS.n1306 AVSS.n1305 585
R416 AVSS.n1405 AVSS.n1404 585
R417 AVSS.n1407 AVSS.n1393 585
R418 AVSS.n1410 AVSS.n1409 585
R419 AVSS.n1391 AVSS.n1390 585
R420 AVSS.n1417 AVSS.n1416 585
R421 AVSS.n1419 AVSS.n1387 585
R422 AVSS.n1422 AVSS.n1421 585
R423 AVSS.n1388 AVSS.n1380 585
R424 AVSS.n1433 AVSS.n1432 585
R425 AVSS.n1435 AVSS.n1379 585
R426 AVSS.n1438 AVSS.n1437 585
R427 AVSS.n1439 AVSS.n1375 585
R428 AVSS.n1446 AVSS.n1445 585
R429 AVSS.n1448 AVSS.n1374 585
R430 AVSS.n1451 AVSS.n1450 585
R431 AVSS.n1452 AVSS.n1370 585
R432 AVSS.n1460 AVSS.n1459 585
R433 AVSS.n1462 AVSS.n1369 585
R434 AVSS.n1463 AVSS.n1362 585
R435 AVSS.n1466 AVSS.n1465 585
R436 AVSS.n1367 AVSS.n1366 585
R437 AVSS.n1365 AVSS.n1355 585
R438 AVSS.n1476 AVSS.n1475 585
R439 AVSS.n1478 AVSS.n1354 585
R440 AVSS.n1481 AVSS.n1480 585
R441 AVSS.n1482 AVSS.n1350 585
R442 AVSS.n1495 AVSS.n1494 585
R443 AVSS.n1497 AVSS.n1349 585
R444 AVSS.n1500 AVSS.n1499 585
R445 AVSS.n1501 AVSS.n1345 585
R446 AVSS.n1509 AVSS.n1508 585
R447 AVSS.n1511 AVSS.n1344 585
R448 AVSS.n1514 AVSS.n1513 585
R449 AVSS.n1341 AVSS.n1340 585
R450 AVSS.n1520 AVSS.n1519 585
R451 AVSS.n1523 AVSS.n1522 585
R452 AVSS.n1339 AVSS.n1335 585
R453 AVSS.n1529 AVSS.n1334 585
R454 AVSS.n1532 AVSS.n1531 585
R455 AVSS.n1534 AVSS.n1331 585
R456 AVSS.n1537 AVSS.n1536 585
R457 AVSS.n1332 AVSS.n1324 585
R458 AVSS.n1547 AVSS.n1546 585
R459 AVSS.n1549 AVSS.n1323 585
R460 AVSS.n1552 AVSS.n1551 585
R461 AVSS.n1320 AVSS.n1319 585
R462 AVSS.n1668 AVSS.n1667 585
R463 AVSS.n1670 AVSS.n1318 585
R464 AVSS.n1673 AVSS.n1672 585
R465 AVSS.n1316 AVSS.n1311 585
R466 AVSS.n1679 AVSS.n1678 585
R467 AVSS.n1680 AVSS.n1679 585
R468 AVSS.n1658 AVSS.n1310 585
R469 AVSS.n1310 AVSS.n1309 585
R470 AVSS.n1657 AVSS.n1656 585
R471 AVSS.n1656 AVSS.n1655 585
R472 AVSS.n1564 AVSS.n1557 585
R473 AVSS.n1558 AVSS.n1557 585
R474 AVSS.n1648 AVSS.n1647 585
R475 AVSS.n1649 AVSS.n1648 585
R476 AVSS.n1563 AVSS.n1562 585
R477 AVSS.n1562 AVSS.n1561 585
R478 AVSS.n1637 AVSS.n1636 585
R479 AVSS.n1636 AVSS.n1290 585
R480 AVSS.n1639 AVSS.n1289 585
R481 AVSS.n1696 AVSS.n1289 585
R482 AVSS.n1635 AVSS.n1288 585
R483 AVSS.n1697 AVSS.n1288 585
R484 AVSS.n1633 AVSS.n1287 585
R485 AVSS.n1698 AVSS.n1287 585
R486 AVSS.n1570 AVSS.n1569 585
R487 AVSS.n1569 AVSS.n1277 585
R488 AVSS.n1628 AVSS.n1276 585
R489 AVSS.n1707 AVSS.n1276 585
R490 AVSS.n1626 AVSS.n1275 585
R491 AVSS.n1708 AVSS.n1275 585
R492 AVSS.n1572 AVSS.n1274 585
R493 AVSS.n1709 AVSS.n1274 585
R494 AVSS.n1620 AVSS.n1619 585
R495 AVSS.n1619 AVSS.n1273 585
R496 AVSS.n1618 AVSS.n1617 585
R497 AVSS.n1618 AVSS.n1255 585
R498 AVSS.n1575 AVSS.n1254 585
R499 AVSS.n1721 AVSS.n1254 585
R500 AVSS.n1597 AVSS.n1253 585
R501 AVSS.n1722 AVSS.n1253 585
R502 AVSS.n1603 AVSS.n1252 585
R503 AVSS.n1723 AVSS.n1252 585
R504 AVSS.n1606 AVSS.n1605 585
R505 AVSS.n1605 AVSS.n1243 585
R506 AVSS.n1595 AVSS.n1242 585
R507 AVSS.n1732 AVSS.n1242 585
R508 AVSS.n1593 AVSS.n1241 585
R509 AVSS.n1733 AVSS.n1241 585
R510 AVSS.n1579 AVSS.n1240 585
R511 AVSS.n1734 AVSS.n1240 585
R512 AVSS.n1588 AVSS.n49 585
R513 AVSS.n51 AVSS.n49 585
R514 AVSS.n1741 AVSS.n50 585
R515 AVSS.n1741 AVSS.n1740 585
R516 AVSS.n1743 AVSS.n1742 585
R517 AVSS.n1742 AVSS.n37 585
R518 AVSS.n48 AVSS.n46 585
R519 AVSS.n48 AVSS.n15 585
R520 AVSS.n1227 AVSS.n1226 585
R521 AVSS.n1228 AVSS.n1227 585
R522 AVSS.n1212 AVSS.n60 585
R523 AVSS.n69 AVSS.n60 585
R524 AVSS.n1211 AVSS.n1210 585
R525 AVSS.n1210 AVSS.n1209 585
R526 AVSS.n1183 AVSS.n67 585
R527 AVSS.n87 AVSS.n67 585
R528 AVSS.n1182 AVSS.n85 585
R529 AVSS.n1192 AVSS.n85 585
R530 AVSS.n105 AVSS.n101 585
R531 AVSS.n107 AVSS.n105 585
R532 AVSS.n1174 AVSS.n1173 585
R533 AVSS.n1173 AVSS.n1172 585
R534 AVSS.n1152 AVSS.n104 585
R535 AVSS.n116 AVSS.n104 585
R536 AVSS.n1151 AVSS.n114 585
R537 AVSS.n1162 AVSS.n114 585
R538 AVSS.n132 AVSS.n126 585
R539 AVSS.n1139 AVSS.n132 585
R540 AVSS.n162 AVSS.n161 585
R541 AVSS.n161 AVSS.n130 585
R542 AVSS.n1066 AVSS.n139 585
R543 AVSS.n1091 AVSS.n139 585
R544 AVSS.n159 AVSS.n158 585
R545 AVSS.n158 AVSS.n157 585
R546 AVSS.n1055 AVSS.n149 585
R547 AVSS.n1074 AVSS.n149 585
R548 AVSS.n1056 AVSS.n1050 585
R549 AVSS.n1050 AVSS.n1049 585
R550 AVSS.n171 AVSS.n170 585
R551 AVSS.n172 AVSS.n171 585
R552 AVSS.n1041 AVSS.n1040 585
R553 AVSS.n1040 AVSS.n1039 585
R554 AVSS.n1018 AVSS.n179 585
R555 AVSS.n195 AVSS.n179 585
R556 AVSS.n1017 AVSS.n193 585
R557 AVSS.n1026 AVSS.n193 585
R558 AVSS.n217 AVSS.n211 585
R559 AVSS.n219 AVSS.n217 585
R560 AVSS.n1007 AVSS.n1006 585
R561 AVSS.n1006 AVSS.n1005 585
R562 AVSS.n216 AVSS.n215 585
R563 AVSS.n234 AVSS.n216 585
R564 AVSS.n986 AVSS.n232 585
R565 AVSS.n993 AVSS.n232 585
R566 AVSS.n984 AVSS.n983 585
R567 AVSS.n983 AVSS.n982 585
R568 AVSS.n970 AVSS.n249 585
R569 AVSS.n250 AVSS.n249 585
R570 AVSS.n969 AVSS.n968 585
R571 AVSS.n968 AVSS.n967 585
R572 AVSS.n259 AVSS.n258 585
R573 AVSS.n279 AVSS.n259 585
R574 AVSS.n912 AVSS.n277 585
R575 AVSS.n933 AVSS.n277 585
R576 AVSS.n914 AVSS.n275 585
R577 AVSS.n945 AVSS.n275 585
R578 AVSS.n289 AVSS.n274 585
R579 AVSS.n946 AVSS.n274 585
R580 AVSS.n922 AVSS.n273 585
R581 AVSS.n947 AVSS.n273 585
R582 AVSS.n745 AVSS.n288 585
R583 AVSS.n746 AVSS.n745 585
R584 AVSS.n744 AVSS.n743 585
R585 AVSS.n753 AVSS.n744 585
R586 AVSS.n329 AVSS.n328 585
R587 AVSS.n754 AVSS.n328 585
R588 AVSS.n737 AVSS.n327 585
R589 AVSS.n755 AVSS.n327 585
R590 AVSS.n735 AVSS.n734 585
R591 AVSS.n734 AVSS.n315 585
R592 AVSS.n331 AVSS.n314 585
R593 AVSS.n765 AVSS.n314 585
R594 AVSS.n728 AVSS.n313 585
R595 AVSS.n766 AVSS.n313 585
R596 AVSS.n333 AVSS.n312 585
R597 AVSS.n767 AVSS.n312 585
R598 AVSS.n721 AVSS.n300 585
R599 AVSS.n302 AVSS.n300 585
R600 AVSS.n779 AVSS.n778 585
R601 AVSS.n778 AVSS.n777 585
R602 AVSS.n299 AVSS.n297 585
R603 AVSS.n301 AVSS.n299 585
R604 AVSS.n715 AVSS.n714 585
R605 AVSS.n714 AVSS.n713 585
R606 AVSS.n339 AVSS.n337 585
R607 AVSS.n340 AVSS.n339 585
R608 AVSS.n699 AVSS.n698 585
R609 AVSS.n700 AVSS.n699 585
R610 AVSS.n697 AVSS.n349 585
R611 AVSS.n349 AVSS.n348 585
R612 AVSS.n354 AVSS.n350 585
R613 AVSS.n356 AVSS.n354 585
R614 AVSS.n692 AVSS.n691 585
R615 AVSS.n691 AVSS.n690 585
R616 AVSS.n379 AVSS.n353 585
R617 AVSS.n355 AVSS.n353 585
R618 AVSS.n674 AVSS.n673 585
R619 AVSS.n675 AVSS.n674 585
R620 AVSS.n661 AVSS.n377 585
R621 AVSS.n680 AVSS.n377 585
R622 AVSS.n663 AVSS.n376 585
R623 AVSS.n681 AVSS.n376 585
R624 AVSS.n660 AVSS.n375 585
R625 AVSS.n682 AVSS.n375 585
R626 AVSS.n391 AVSS.n382 585
R627 AVSS.n391 AVSS.n374 585
R628 AVSS.n652 AVSS.n651 585
R629 AVSS.n651 AVSS.n650 585
R630 AVSS.n390 AVSS.n387 585
R631 AVSS.n392 AVSS.n390 585
R632 AVSS.n516 AVSS.n515 585
R633 AVSS.n518 AVSS.n508 585
R634 AVSS.n520 AVSS.n519 585
R635 AVSS.n502 AVSS.n500 585
R636 AVSS.n531 AVSS.n530 585
R637 AVSS.n533 AVSS.n498 585
R638 AVSS.n535 AVSS.n534 585
R639 AVSS.n495 AVSS.n493 585
R640 AVSS.n542 AVSS.n541 585
R641 AVSS.n544 AVSS.n492 585
R642 AVSS.n546 AVSS.n545 585
R643 AVSS.n487 AVSS.n485 585
R644 AVSS.n552 AVSS.n551 585
R645 AVSS.n554 AVSS.n484 585
R646 AVSS.n556 AVSS.n555 585
R647 AVSS.n472 AVSS.n470 585
R648 AVSS.n563 AVSS.n562 585
R649 AVSS.n565 AVSS.n469 585
R650 AVSS.n567 AVSS.n566 585
R651 AVSS.n464 AVSS.n462 585
R652 AVSS.n573 AVSS.n572 585
R653 AVSS.n575 AVSS.n461 585
R654 AVSS.n577 AVSS.n576 585
R655 AVSS.n459 AVSS.n453 585
R656 AVSS.n458 AVSS.n457 585
R657 AVSS.n444 AVSS.n442 585
R658 AVSS.n586 AVSS.n585 585
R659 AVSS.n588 AVSS.n441 585
R660 AVSS.n590 AVSS.n589 585
R661 AVSS.n436 AVSS.n434 585
R662 AVSS.n596 AVSS.n595 585
R663 AVSS.n598 AVSS.n433 585
R664 AVSS.n600 AVSS.n599 585
R665 AVSS.n427 AVSS.n425 585
R666 AVSS.n606 AVSS.n605 585
R667 AVSS.n608 AVSS.n424 585
R668 AVSS.n610 AVSS.n609 585
R669 AVSS.n418 AVSS.n417 585
R670 AVSS.n621 AVSS.n620 585
R671 AVSS.n624 AVSS.n623 585
R672 AVSS.n416 AVSS.n411 585
R673 AVSS.n629 AVSS.n409 585
R674 AVSS.n631 AVSS.n630 585
R675 AVSS.n633 AVSS.n404 585
R676 AVSS.n635 AVSS.n634 585
R677 AVSS.n405 AVSS.n401 585
R678 AVSS.n406 AVSS.n394 585
R679 AVSS.n643 AVSS.n393 585
R680 AVSS.n647 AVSS.n646 585
R681 AVSS.n647 AVSS.n392 585
R682 AVSS.n649 AVSS.n648 585
R683 AVSS.n650 AVSS.n649 585
R684 AVSS.n371 AVSS.n370 585
R685 AVSS.n374 AVSS.n371 585
R686 AVSS.n684 AVSS.n683 585
R687 AVSS.n683 AVSS.n682 585
R688 AVSS.n373 AVSS.n372 585
R689 AVSS.n681 AVSS.n373 585
R690 AVSS.n679 AVSS.n678 585
R691 AVSS.n680 AVSS.n679 585
R692 AVSS.n677 AVSS.n676 585
R693 AVSS.n677 AVSS.n675 585
R694 AVSS.n364 AVSS.n357 585
R695 AVSS.n357 AVSS.n355 585
R696 AVSS.n689 AVSS.n688 585
R697 AVSS.n690 AVSS.n689 585
R698 AVSS.n360 AVSS.n358 585
R699 AVSS.n358 AVSS.n356 585
R700 AVSS.n347 AVSS.n345 585
R701 AVSS.n348 AVSS.n347 585
R702 AVSS.n702 AVSS.n701 585
R703 AVSS.n701 AVSS.n700 585
R704 AVSS.n346 AVSS.n341 585
R705 AVSS.n341 AVSS.n340 585
R706 AVSS.n712 AVSS.n711 585
R707 AVSS.n713 AVSS.n712 585
R708 AVSS.n343 AVSS.n303 585
R709 AVSS.n303 AVSS.n301 585
R710 AVSS.n776 AVSS.n775 585
R711 AVSS.n777 AVSS.n776 585
R712 AVSS.n306 AVSS.n304 585
R713 AVSS.n304 AVSS.n302 585
R714 AVSS.n769 AVSS.n768 585
R715 AVSS.n768 AVSS.n767 585
R716 AVSS.n317 AVSS.n311 585
R717 AVSS.n766 AVSS.n311 585
R718 AVSS.n764 AVSS.n763 585
R719 AVSS.n765 AVSS.n764 585
R720 AVSS.n319 AVSS.n316 585
R721 AVSS.n316 AVSS.n315 585
R722 AVSS.n757 AVSS.n756 585
R723 AVSS.n756 AVSS.n755 585
R724 AVSS.n747 AVSS.n326 585
R725 AVSS.n754 AVSS.n326 585
R726 AVSS.n752 AVSS.n751 585
R727 AVSS.n753 AVSS.n752 585
R728 AVSS.n270 AVSS.n268 585
R729 AVSS.n746 AVSS.n270 585
R730 AVSS.n949 AVSS.n948 585
R731 AVSS.n948 AVSS.n947 585
R732 AVSS.n935 AVSS.n271 585
R733 AVSS.n946 AVSS.n271 585
R734 AVSS.n944 AVSS.n943 585
R735 AVSS.n945 AVSS.n944 585
R736 AVSS.n941 AVSS.n934 585
R737 AVSS.n934 AVSS.n933 585
R738 AVSS.n263 AVSS.n261 585
R739 AVSS.n279 AVSS.n261 585
R740 AVSS.n966 AVSS.n965 585
R741 AVSS.n967 AVSS.n966 585
R742 AVSS.n264 AVSS.n262 585
R743 AVSS.n262 AVSS.n250 585
R744 AVSS.n958 AVSS.n230 585
R745 AVSS.n982 AVSS.n230 585
R746 AVSS.n995 AVSS.n994 585
R747 AVSS.n994 AVSS.n993 585
R748 AVSS.n996 AVSS.n221 585
R749 AVSS.n234 AVSS.n221 585
R750 AVSS.n1004 AVSS.n1003 585
R751 AVSS.n1005 AVSS.n1004 585
R752 AVSS.n223 AVSS.n191 585
R753 AVSS.n219 AVSS.n191 585
R754 AVSS.n1028 AVSS.n1027 585
R755 AVSS.n1027 AVSS.n1026 585
R756 AVSS.n1029 AVSS.n181 585
R757 AVSS.n195 AVSS.n181 585
R758 AVSS.n1038 AVSS.n1037 585
R759 AVSS.n1039 AVSS.n1038 585
R760 AVSS.n184 AVSS.n182 585
R761 AVSS.n182 AVSS.n172 585
R762 AVSS.n147 AVSS.n146 585
R763 AVSS.n1049 AVSS.n147 585
R764 AVSS.n1076 AVSS.n1075 585
R765 AVSS.n1075 AVSS.n1074 585
R766 AVSS.n1077 AVSS.n140 585
R767 AVSS.n157 AVSS.n140 585
R768 AVSS.n1090 AVSS.n1089 585
R769 AVSS.n1091 AVSS.n1090 585
R770 AVSS.n143 AVSS.n141 585
R771 AVSS.n141 AVSS.n130 585
R772 AVSS.n1083 AVSS.n113 585
R773 AVSS.n1139 AVSS.n113 585
R774 AVSS.n1164 AVSS.n1163 585
R775 AVSS.n1163 AVSS.n1162 585
R776 AVSS.n110 AVSS.n109 585
R777 AVSS.n116 AVSS.n109 585
R778 AVSS.n1171 AVSS.n1170 585
R779 AVSS.n1172 AVSS.n1171 585
R780 AVSS.n83 AVSS.n77 585
R781 AVSS.n107 AVSS.n83 585
R782 AVSS.n1194 AVSS.n1193 585
R783 AVSS.n1193 AVSS.n1192 585
R784 AVSS.n78 AVSS.n71 585
R785 AVSS.n87 AVSS.n71 585
R786 AVSS.n1208 AVSS.n1207 585
R787 AVSS.n1209 AVSS.n1208 585
R788 AVSS.n73 AVSS.n57 585
R789 AVSS.n69 AVSS.n57 585
R790 AVSS.n1229 AVSS.n58 585
R791 AVSS.n1229 AVSS.n1228 585
R792 AVSS.n1231 AVSS.n1230 585
R793 AVSS.n1230 AVSS.n15 585
R794 AVSS.n1232 AVSS.n52 585
R795 AVSS.n52 AVSS.n37 585
R796 AVSS.n1739 AVSS.n1738 585
R797 AVSS.n1740 AVSS.n1739 585
R798 AVSS.n1737 AVSS.n53 585
R799 AVSS.n53 AVSS.n51 585
R800 AVSS.n1736 AVSS.n1735 585
R801 AVSS.n1735 AVSS.n1734 585
R802 AVSS.n1245 AVSS.n1239 585
R803 AVSS.n1733 AVSS.n1239 585
R804 AVSS.n1731 AVSS.n1730 585
R805 AVSS.n1732 AVSS.n1731 585
R806 AVSS.n1247 AVSS.n1244 585
R807 AVSS.n1244 AVSS.n1243 585
R808 AVSS.n1725 AVSS.n1724 585
R809 AVSS.n1724 AVSS.n1723 585
R810 AVSS.n1257 AVSS.n1251 585
R811 AVSS.n1722 AVSS.n1251 585
R812 AVSS.n1720 AVSS.n1719 585
R813 AVSS.n1721 AVSS.n1720 585
R814 AVSS.n1259 AVSS.n1256 585
R815 AVSS.n1256 AVSS.n1255 585
R816 AVSS.n1271 AVSS.n1269 585
R817 AVSS.n1273 AVSS.n1271 585
R818 AVSS.n1711 AVSS.n1710 585
R819 AVSS.n1710 AVSS.n1709 585
R820 AVSS.n1279 AVSS.n1272 585
R821 AVSS.n1708 AVSS.n1272 585
R822 AVSS.n1706 AVSS.n1705 585
R823 AVSS.n1707 AVSS.n1706 585
R824 AVSS.n1281 AVSS.n1278 585
R825 AVSS.n1278 AVSS.n1277 585
R826 AVSS.n1700 AVSS.n1699 585
R827 AVSS.n1699 AVSS.n1698 585
R828 AVSS.n1292 AVSS.n1286 585
R829 AVSS.n1697 AVSS.n1286 585
R830 AVSS.n1695 AVSS.n1694 585
R831 AVSS.n1696 AVSS.n1695 585
R832 AVSS.n1294 AVSS.n1291 585
R833 AVSS.n1291 AVSS.n1290 585
R834 AVSS.n1559 AVSS.n1297 585
R835 AVSS.n1561 AVSS.n1559 585
R836 AVSS.n1650 AVSS.n1560 585
R837 AVSS.n1650 AVSS.n1649 585
R838 AVSS.n1652 AVSS.n1651 585
R839 AVSS.n1652 AVSS.n1558 585
R840 AVSS.n1654 AVSS.n1653 585
R841 AVSS.n1655 AVSS.n1654 585
R842 AVSS.n1308 AVSS.n1307 585
R843 AVSS.n1309 AVSS.n1308 585
R844 AVSS.n1681 AVSS.n1301 585
R845 AVSS.n1681 AVSS.n1680 585
R846 AVSS.n873 AVSS.n872 585
R847 AVSS.n876 AVSS.n875 585
R848 AVSS.n878 AVSS.n877 585
R849 AVSS.n881 AVSS.n880 585
R850 AVSS.n883 AVSS.n882 585
R851 AVSS.n886 AVSS.n885 585
R852 AVSS.n897 AVSS.n896 585
R853 AVSS.n894 AVSS.n792 585
R854 AVSS.n893 AVSS.n887 585
R855 AVSS.n891 AVSS.n890 585
R856 AVSS.n889 AVSS.n293 585
R857 AVSS.n901 AVSS.n292 585
R858 AVSS.n904 AVSS.n903 585
R859 AVSS.n907 AVSS.n906 585
R860 AVSS.n909 AVSS.n280 585
R861 AVSS.n280 AVSS.n276 585
R862 AVSS.n931 AVSS.n930 585
R863 AVSS.n932 AVSS.n931 585
R864 AVSS.n283 AVSS.n281 585
R865 AVSS.n281 AVSS.n260 585
R866 AVSS.n253 AVSS.n252 585
R867 AVSS.t52 AVSS.n252 585
R868 AVSS.n980 AVSS.n979 585
R869 AVSS.n981 AVSS.n980 585
R870 AVSS.n254 AVSS.n235 585
R871 AVSS.n235 AVSS.n231 585
R872 AVSS.n991 AVSS.n990 585
R873 AVSS.n992 AVSS.n991 585
R874 AVSS.n238 AVSS.n236 585
R875 AVSS.n236 AVSS.n218 585
R876 AVSS.n244 AVSS.n243 585
R877 AVSS.n243 AVSS.n220 585
R878 AVSS.n241 AVSS.n196 585
R879 AVSS.n196 AVSS.n192 585
R880 AVSS.n1024 AVSS.n1023 585
R881 AVSS.n1025 AVSS.n1024 585
R882 AVSS.n199 AVSS.n197 585
R883 AVSS.n812 AVSS.n197 585
R884 AVSS.n202 AVSS.n174 585
R885 AVSS.n180 AVSS.n174 585
R886 AVSS.n1047 AVSS.n1046 585
R887 AVSS.n1048 AVSS.n1047 585
R888 AVSS.n176 AVSS.n151 585
R889 AVSS.n151 AVSS.n148 585
R890 AVSS.n1072 AVSS.n1071 585
R891 AVSS.n1073 AVSS.n1072 585
R892 AVSS.n154 AVSS.n152 585
R893 AVSS.n152 AVSS.n138 585
R894 AVSS.n165 AVSS.n129 585
R895 AVSS.n1092 AVSS.n129 585
R896 AVSS.n1142 AVSS.n1141 585
R897 AVSS.n1141 AVSS.n1140 585
R898 AVSS.n1143 AVSS.n117 585
R899 AVSS.n1138 AVSS.n117 585
R900 AVSS.n1160 AVSS.n1159 585
R901 AVSS.n1161 AVSS.n1160 585
R902 AVSS.n124 AVSS.n118 585
R903 AVSS.n118 AVSS.n106 585
R904 AVSS.n123 AVSS.n122 585
R905 AVSS.n122 AVSS.n108 585
R906 AVSS.n120 AVSS.n88 585
R907 AVSS.n88 AVSS.n84 585
R908 AVSS.n1190 AVSS.n1189 585
R909 AVSS.n1191 AVSS.n1190 585
R910 AVSS.n92 AVSS.n90 585
R911 AVSS.n90 AVSS.n68 585
R912 AVSS.n89 AVSS.n64 585
R913 AVSS.n89 AVSS.n70 585
R914 AVSS.n1217 AVSS.n42 585
R915 AVSS.n59 AVSS.n42 585
R916 AVSS.n1751 AVSS.n1750 585
R917 AVSS.n44 AVSS.n41 585
R918 AVSS.n1746 AVSS.n40 585
R919 AVSS.n1753 AVSS.n40 585
R920 AVSS.n39 AVSS.n38 585
R921 AVSS.n19 AVSS.n18 585
R922 AVSS.n21 AVSS.n20 585
R923 AVSS.n23 AVSS.n22 585
R924 AVSS.n25 AVSS.n24 585
R925 AVSS.n28 AVSS.n27 585
R926 AVSS.n30 AVSS.n29 585
R927 AVSS.n33 AVSS.n32 585
R928 AVSS.n35 AVSS.n34 585
R929 AVSS.n13 AVSS.n11 585
R930 AVSS.n1755 AVSS.n1754 585
R931 AVSS.n1754 AVSS.n1753 585
R932 AVSS.n1108 AVSS.n14 585
R933 AVSS.n59 AVSS.n14 585
R934 AVSS.n1118 AVSS.n1117 585
R935 AVSS.n1118 AVSS.n70 585
R936 AVSS.n1120 AVSS.n1119 585
R937 AVSS.n1119 AVSS.n68 585
R938 AVSS.n1103 AVSS.n86 585
R939 AVSS.n1191 AVSS.n86 585
R940 AVSS.n1126 AVSS.n1125 585
R941 AVSS.n1126 AVSS.n84 585
R942 AVSS.n1127 AVSS.n1101 585
R943 AVSS.n1127 AVSS.n108 585
R944 AVSS.n1129 AVSS.n1128 585
R945 AVSS.n1128 AVSS.n106 585
R946 AVSS.n134 AVSS.n115 585
R947 AVSS.n1161 AVSS.n115 585
R948 AVSS.n1137 AVSS.n1136 585
R949 AVSS.n1138 AVSS.n1137 585
R950 AVSS.n1095 AVSS.n131 585
R951 AVSS.n1140 AVSS.n131 585
R952 AVSS.n1094 AVSS.n1093 585
R953 AVSS.n1093 AVSS.n1092 585
R954 AVSS.n823 AVSS.n137 585
R955 AVSS.n138 AVSS.n137 585
R956 AVSS.n816 AVSS.n150 585
R957 AVSS.n1073 AVSS.n150 585
R958 AVSS.n833 AVSS.n832 585
R959 AVSS.n832 AVSS.n148 585
R960 AVSS.n835 AVSS.n173 585
R961 AVSS.n1048 AVSS.n173 585
R962 AVSS.n815 AVSS.n814 585
R963 AVSS.n814 AVSS.n180 585
R964 AVSS.n813 AVSS.n808 585
R965 AVSS.n813 AVSS.n812 585
R966 AVSS.n843 AVSS.n194 585
R967 AVSS.n1025 AVSS.n194 585
R968 AVSS.n805 AVSS.n804 585
R969 AVSS.n804 AVSS.n192 585
R970 AVSS.n851 AVSS.n850 585
R971 AVSS.n851 AVSS.n220 585
R972 AVSS.n853 AVSS.n852 585
R973 AVSS.n852 AVSS.n218 585
R974 AVSS.n855 AVSS.n233 585
R975 AVSS.n992 AVSS.n233 585
R976 AVSS.n801 AVSS.n800 585
R977 AVSS.n800 AVSS.n231 585
R978 AVSS.n860 AVSS.n251 585
R979 AVSS.n981 AVSS.n251 585
R980 AVSS.n863 AVSS.n862 585
R981 AVSS.n862 AVSS.t52 585
R982 AVSS.n861 AVSS.n799 585
R983 AVSS.n861 AVSS.n260 585
R984 AVSS.n794 AVSS.n278 585
R985 AVSS.n932 AVSS.n278 585
R986 AVSS.n871 AVSS.n793 585
R987 AVSS.n793 AVSS.n276 585
R988 AVSS.n891 AVSS.n889 538.854
R989 AVSS.n649 AVSS.n647 394
R990 AVSS.n649 AVSS.n371 394
R991 AVSS.n683 AVSS.n371 394
R992 AVSS.n683 AVSS.n373 394
R993 AVSS.n679 AVSS.n373 394
R994 AVSS.n679 AVSS.n677 394
R995 AVSS.n677 AVSS.n357 394
R996 AVSS.n689 AVSS.n357 394
R997 AVSS.n689 AVSS.n358 394
R998 AVSS.n358 AVSS.n347 394
R999 AVSS.n701 AVSS.n347 394
R1000 AVSS.n701 AVSS.n341 394
R1001 AVSS.n712 AVSS.n341 394
R1002 AVSS.n712 AVSS.n303 394
R1003 AVSS.n776 AVSS.n303 394
R1004 AVSS.n776 AVSS.n304 394
R1005 AVSS.n768 AVSS.n304 394
R1006 AVSS.n768 AVSS.n311 394
R1007 AVSS.n764 AVSS.n311 394
R1008 AVSS.n764 AVSS.n316 394
R1009 AVSS.n756 AVSS.n316 394
R1010 AVSS.n756 AVSS.n326 394
R1011 AVSS.n752 AVSS.n326 394
R1012 AVSS.n752 AVSS.n270 394
R1013 AVSS.n948 AVSS.n270 394
R1014 AVSS.n948 AVSS.n271 394
R1015 AVSS.n944 AVSS.n271 394
R1016 AVSS.n944 AVSS.n934 394
R1017 AVSS.n934 AVSS.n261 394
R1018 AVSS.n966 AVSS.n261 394
R1019 AVSS.n966 AVSS.n262 394
R1020 AVSS.n262 AVSS.n230 394
R1021 AVSS.n994 AVSS.n230 394
R1022 AVSS.n994 AVSS.n221 394
R1023 AVSS.n1004 AVSS.n221 394
R1024 AVSS.n1004 AVSS.n191 394
R1025 AVSS.n1027 AVSS.n191 394
R1026 AVSS.n1027 AVSS.n181 394
R1027 AVSS.n1038 AVSS.n181 394
R1028 AVSS.n1038 AVSS.n182 394
R1029 AVSS.n182 AVSS.n147 394
R1030 AVSS.n1075 AVSS.n147 394
R1031 AVSS.n1075 AVSS.n140 394
R1032 AVSS.n1090 AVSS.n140 394
R1033 AVSS.n1090 AVSS.n141 394
R1034 AVSS.n141 AVSS.n113 394
R1035 AVSS.n1163 AVSS.n113 394
R1036 AVSS.n1163 AVSS.n109 394
R1037 AVSS.n1171 AVSS.n109 394
R1038 AVSS.n1171 AVSS.n83 394
R1039 AVSS.n1193 AVSS.n83 394
R1040 AVSS.n1193 AVSS.n71 394
R1041 AVSS.n1208 AVSS.n71 394
R1042 AVSS.n1208 AVSS.n57 394
R1043 AVSS.n1229 AVSS.n57 394
R1044 AVSS.n1230 AVSS.n1229 394
R1045 AVSS.n1230 AVSS.n52 394
R1046 AVSS.n1739 AVSS.n52 394
R1047 AVSS.n1739 AVSS.n53 394
R1048 AVSS.n1735 AVSS.n53 394
R1049 AVSS.n1735 AVSS.n1239 394
R1050 AVSS.n1731 AVSS.n1239 394
R1051 AVSS.n1731 AVSS.n1244 394
R1052 AVSS.n1724 AVSS.n1244 394
R1053 AVSS.n1724 AVSS.n1251 394
R1054 AVSS.n1720 AVSS.n1251 394
R1055 AVSS.n1720 AVSS.n1256 394
R1056 AVSS.n1271 AVSS.n1256 394
R1057 AVSS.n1710 AVSS.n1271 394
R1058 AVSS.n1710 AVSS.n1272 394
R1059 AVSS.n1706 AVSS.n1272 394
R1060 AVSS.n1706 AVSS.n1278 394
R1061 AVSS.n1699 AVSS.n1278 394
R1062 AVSS.n1699 AVSS.n1286 394
R1063 AVSS.n1695 AVSS.n1286 394
R1064 AVSS.n1695 AVSS.n1291 394
R1065 AVSS.n1559 AVSS.n1291 394
R1066 AVSS.n1650 AVSS.n1559 394
R1067 AVSS.n1652 AVSS.n1650 394
R1068 AVSS.n1654 AVSS.n1652 394
R1069 AVSS.n1654 AVSS.n1308 394
R1070 AVSS.n1681 AVSS.n1308 394
R1071 AVSS.n406 AVSS.n405 394
R1072 AVSS.n634 AVSS.n633 394
R1073 AVSS.n631 AVSS.n409 394
R1074 AVSS.n623 AVSS.n416 394
R1075 AVSS.n621 AVSS.n417 394
R1076 AVSS.n609 AVSS.n608 394
R1077 AVSS.n606 AVSS.n425 394
R1078 AVSS.n599 AVSS.n598 394
R1079 AVSS.n596 AVSS.n434 394
R1080 AVSS.n589 AVSS.n588 394
R1081 AVSS.n586 AVSS.n442 394
R1082 AVSS.n459 AVSS.n458 394
R1083 AVSS.n576 AVSS.n575 394
R1084 AVSS.n573 AVSS.n462 394
R1085 AVSS.n566 AVSS.n565 394
R1086 AVSS.n563 AVSS.n470 394
R1087 AVSS.n555 AVSS.n554 394
R1088 AVSS.n552 AVSS.n485 394
R1089 AVSS.n545 AVSS.n544 394
R1090 AVSS.n542 AVSS.n493 394
R1091 AVSS.n534 AVSS.n533 394
R1092 AVSS.n531 AVSS.n500 394
R1093 AVSS.n519 AVSS.n518 394
R1094 AVSS.n651 AVSS.n390 394
R1095 AVSS.n651 AVSS.n391 394
R1096 AVSS.n391 AVSS.n375 394
R1097 AVSS.n376 AVSS.n375 394
R1098 AVSS.n377 AVSS.n376 394
R1099 AVSS.n674 AVSS.n377 394
R1100 AVSS.n674 AVSS.n353 394
R1101 AVSS.n691 AVSS.n353 394
R1102 AVSS.n691 AVSS.n354 394
R1103 AVSS.n354 AVSS.n349 394
R1104 AVSS.n699 AVSS.n349 394
R1105 AVSS.n699 AVSS.n339 394
R1106 AVSS.n714 AVSS.n339 394
R1107 AVSS.n714 AVSS.n299 394
R1108 AVSS.n778 AVSS.n299 394
R1109 AVSS.n778 AVSS.n300 394
R1110 AVSS.n312 AVSS.n300 394
R1111 AVSS.n313 AVSS.n312 394
R1112 AVSS.n314 AVSS.n313 394
R1113 AVSS.n734 AVSS.n314 394
R1114 AVSS.n734 AVSS.n327 394
R1115 AVSS.n328 AVSS.n327 394
R1116 AVSS.n744 AVSS.n328 394
R1117 AVSS.n745 AVSS.n744 394
R1118 AVSS.n745 AVSS.n273 394
R1119 AVSS.n274 AVSS.n273 394
R1120 AVSS.n275 AVSS.n274 394
R1121 AVSS.n277 AVSS.n275 394
R1122 AVSS.n277 AVSS.n259 394
R1123 AVSS.n968 AVSS.n259 394
R1124 AVSS.n968 AVSS.n249 394
R1125 AVSS.n983 AVSS.n249 394
R1126 AVSS.n983 AVSS.n232 394
R1127 AVSS.n232 AVSS.n216 394
R1128 AVSS.n1006 AVSS.n216 394
R1129 AVSS.n1006 AVSS.n217 394
R1130 AVSS.n217 AVSS.n193 394
R1131 AVSS.n193 AVSS.n179 394
R1132 AVSS.n1040 AVSS.n179 394
R1133 AVSS.n1040 AVSS.n171 394
R1134 AVSS.n1050 AVSS.n171 394
R1135 AVSS.n1050 AVSS.n149 394
R1136 AVSS.n158 AVSS.n149 394
R1137 AVSS.n158 AVSS.n139 394
R1138 AVSS.n161 AVSS.n139 394
R1139 AVSS.n161 AVSS.n132 394
R1140 AVSS.n132 AVSS.n114 394
R1141 AVSS.n114 AVSS.n104 394
R1142 AVSS.n1173 AVSS.n104 394
R1143 AVSS.n1173 AVSS.n105 394
R1144 AVSS.n105 AVSS.n85 394
R1145 AVSS.n85 AVSS.n67 394
R1146 AVSS.n1210 AVSS.n67 394
R1147 AVSS.n1210 AVSS.n60 394
R1148 AVSS.n1227 AVSS.n60 394
R1149 AVSS.n1227 AVSS.n48 394
R1150 AVSS.n1742 AVSS.n48 394
R1151 AVSS.n1742 AVSS.n1741 394
R1152 AVSS.n1741 AVSS.n49 394
R1153 AVSS.n1240 AVSS.n49 394
R1154 AVSS.n1241 AVSS.n1240 394
R1155 AVSS.n1242 AVSS.n1241 394
R1156 AVSS.n1605 AVSS.n1242 394
R1157 AVSS.n1605 AVSS.n1252 394
R1158 AVSS.n1253 AVSS.n1252 394
R1159 AVSS.n1254 AVSS.n1253 394
R1160 AVSS.n1618 AVSS.n1254 394
R1161 AVSS.n1619 AVSS.n1618 394
R1162 AVSS.n1619 AVSS.n1274 394
R1163 AVSS.n1275 AVSS.n1274 394
R1164 AVSS.n1276 AVSS.n1275 394
R1165 AVSS.n1569 AVSS.n1276 394
R1166 AVSS.n1569 AVSS.n1287 394
R1167 AVSS.n1288 AVSS.n1287 394
R1168 AVSS.n1289 AVSS.n1288 394
R1169 AVSS.n1636 AVSS.n1289 394
R1170 AVSS.n1636 AVSS.n1562 394
R1171 AVSS.n1648 AVSS.n1562 394
R1172 AVSS.n1648 AVSS.n1557 394
R1173 AVSS.n1656 AVSS.n1557 394
R1174 AVSS.n1656 AVSS.n1310 394
R1175 AVSS.n1679 AVSS.n1310 394
R1176 AVSS.n1684 AVSS.n1305 394
R1177 AVSS.n1405 AVSS.n1305 394
R1178 AVSS.n1409 AVSS.n1407 394
R1179 AVSS.n1417 AVSS.n1390 394
R1180 AVSS.n1421 AVSS.n1419 394
R1181 AVSS.n1433 AVSS.n1380 394
R1182 AVSS.n1437 AVSS.n1435 394
R1183 AVSS.n1446 AVSS.n1375 394
R1184 AVSS.n1450 AVSS.n1448 394
R1185 AVSS.n1460 AVSS.n1370 394
R1186 AVSS.n1463 AVSS.n1462 394
R1187 AVSS.n1465 AVSS.n1367 394
R1188 AVSS.n1476 AVSS.n1355 394
R1189 AVSS.n1480 AVSS.n1478 394
R1190 AVSS.n1495 AVSS.n1350 394
R1191 AVSS.n1499 AVSS.n1497 394
R1192 AVSS.n1509 AVSS.n1345 394
R1193 AVSS.n1513 AVSS.n1511 394
R1194 AVSS.n1520 AVSS.n1340 394
R1195 AVSS.n1522 AVSS.n1339 394
R1196 AVSS.n1532 AVSS.n1334 394
R1197 AVSS.n1536 AVSS.n1534 394
R1198 AVSS.n1547 AVSS.n1324 394
R1199 AVSS.n1551 AVSS.n1549 394
R1200 AVSS.n1668 AVSS.n1319 394
R1201 AVSS.n1672 AVSS.n1670 394
R1202 AVSS.n931 AVSS.n280 394
R1203 AVSS.n931 AVSS.n281 394
R1204 AVSS.n281 AVSS.n252 394
R1205 AVSS.n980 AVSS.n252 394
R1206 AVSS.n980 AVSS.n235 394
R1207 AVSS.n991 AVSS.n235 394
R1208 AVSS.n991 AVSS.n236 394
R1209 AVSS.n243 AVSS.n236 394
R1210 AVSS.n243 AVSS.n196 394
R1211 AVSS.n1024 AVSS.n196 394
R1212 AVSS.n1024 AVSS.n197 394
R1213 AVSS.n197 AVSS.n174 394
R1214 AVSS.n1047 AVSS.n174 394
R1215 AVSS.n1047 AVSS.n151 394
R1216 AVSS.n1072 AVSS.n151 394
R1217 AVSS.n1072 AVSS.n152 394
R1218 AVSS.n152 AVSS.n129 394
R1219 AVSS.n1141 AVSS.n129 394
R1220 AVSS.n1141 AVSS.n117 394
R1221 AVSS.n1160 AVSS.n117 394
R1222 AVSS.n1160 AVSS.n118 394
R1223 AVSS.n122 AVSS.n118 394
R1224 AVSS.n122 AVSS.n88 394
R1225 AVSS.n1190 AVSS.n88 394
R1226 AVSS.n1190 AVSS.n90 394
R1227 AVSS.n90 AVSS.n89 394
R1228 AVSS.n89 AVSS.n42 394
R1229 AVSS.n41 AVSS.n40 394
R1230 AVSS.n40 AVSS.n39 394
R1231 AVSS.n20 AVSS.n19 394
R1232 AVSS.n25 AVSS.n23 394
R1233 AVSS.n30 AVSS.n28 394
R1234 AVSS.n35 AVSS.n33 394
R1235 AVSS.n1754 AVSS.n13 394
R1236 AVSS.n793 AVSS.n278 394
R1237 AVSS.n861 AVSS.n278 394
R1238 AVSS.n862 AVSS.n861 394
R1239 AVSS.n862 AVSS.n251 394
R1240 AVSS.n800 AVSS.n251 394
R1241 AVSS.n800 AVSS.n233 394
R1242 AVSS.n852 AVSS.n233 394
R1243 AVSS.n852 AVSS.n851 394
R1244 AVSS.n851 AVSS.n804 394
R1245 AVSS.n804 AVSS.n194 394
R1246 AVSS.n813 AVSS.n194 394
R1247 AVSS.n814 AVSS.n813 394
R1248 AVSS.n814 AVSS.n173 394
R1249 AVSS.n832 AVSS.n173 394
R1250 AVSS.n832 AVSS.n150 394
R1251 AVSS.n150 AVSS.n137 394
R1252 AVSS.n1093 AVSS.n137 394
R1253 AVSS.n1093 AVSS.n131 394
R1254 AVSS.n1137 AVSS.n131 394
R1255 AVSS.n1137 AVSS.n115 394
R1256 AVSS.n1128 AVSS.n115 394
R1257 AVSS.n1128 AVSS.n1127 394
R1258 AVSS.n1127 AVSS.n1126 394
R1259 AVSS.n1126 AVSS.n86 394
R1260 AVSS.n1119 AVSS.n86 394
R1261 AVSS.n1119 AVSS.n1118 394
R1262 AVSS.n1118 AVSS.n14 394
R1263 AVSS.n904 AVSS.n292 394
R1264 AVSS.n894 AVSS.n893 394
R1265 AVSS.n896 AVSS.n886 394
R1266 AVSS.n883 AVSS.n881 394
R1267 AVSS.n878 AVSS.n876 394
R1268 AVSS.n1683 AVSS.n1306 218.815
R1269 AVSS.n1406 AVSS.n1306 218.815
R1270 AVSS.n1408 AVSS.n1306 218.815
R1271 AVSS.n1418 AVSS.n1306 218.815
R1272 AVSS.n1420 AVSS.n1306 218.815
R1273 AVSS.n1434 AVSS.n1306 218.815
R1274 AVSS.n1436 AVSS.n1306 218.815
R1275 AVSS.n1447 AVSS.n1306 218.815
R1276 AVSS.n1449 AVSS.n1306 218.815
R1277 AVSS.n1461 AVSS.n1306 218.815
R1278 AVSS.n1464 AVSS.n1306 218.815
R1279 AVSS.n1364 AVSS.n1306 218.815
R1280 AVSS.n1477 AVSS.n1306 218.815
R1281 AVSS.n1479 AVSS.n1306 218.815
R1282 AVSS.n1496 AVSS.n1306 218.815
R1283 AVSS.n1498 AVSS.n1306 218.815
R1284 AVSS.n1510 AVSS.n1306 218.815
R1285 AVSS.n1512 AVSS.n1306 218.815
R1286 AVSS.n1521 AVSS.n1306 218.815
R1287 AVSS.n1338 AVSS.n1306 218.815
R1288 AVSS.n1533 AVSS.n1306 218.815
R1289 AVSS.n1535 AVSS.n1306 218.815
R1290 AVSS.n1548 AVSS.n1306 218.815
R1291 AVSS.n1550 AVSS.n1306 218.815
R1292 AVSS.n1669 AVSS.n1306 218.815
R1293 AVSS.n1671 AVSS.n1306 218.815
R1294 AVSS.n517 AVSS.n408 218.815
R1295 AVSS.n507 AVSS.n408 218.815
R1296 AVSS.n532 AVSS.n408 218.815
R1297 AVSS.n499 AVSS.n408 218.815
R1298 AVSS.n543 AVSS.n408 218.815
R1299 AVSS.n491 AVSS.n408 218.815
R1300 AVSS.n553 AVSS.n408 218.815
R1301 AVSS.n483 AVSS.n408 218.815
R1302 AVSS.n564 AVSS.n408 218.815
R1303 AVSS.n468 AVSS.n408 218.815
R1304 AVSS.n574 AVSS.n408 218.815
R1305 AVSS.n460 AVSS.n408 218.815
R1306 AVSS.n455 AVSS.n408 218.815
R1307 AVSS.n587 AVSS.n408 218.815
R1308 AVSS.n440 AVSS.n408 218.815
R1309 AVSS.n597 AVSS.n408 218.815
R1310 AVSS.n432 AVSS.n408 218.815
R1311 AVSS.n607 AVSS.n408 218.815
R1312 AVSS.n423 AVSS.n408 218.815
R1313 AVSS.n622 AVSS.n408 218.815
R1314 AVSS.n415 AVSS.n408 218.815
R1315 AVSS.n632 AVSS.n408 218.815
R1316 AVSS.n408 AVSS.n403 218.815
R1317 AVSS.n408 AVSS.n407 218.815
R1318 AVSS.n874 AVSS.n272 218.815
R1319 AVSS.n879 AVSS.n272 218.815
R1320 AVSS.n884 AVSS.n272 218.815
R1321 AVSS.n895 AVSS.n272 218.815
R1322 AVSS.n892 AVSS.n272 218.815
R1323 AVSS.n888 AVSS.n272 218.815
R1324 AVSS.n905 AVSS.n272 218.815
R1325 AVSS.n1753 AVSS.n1752 218.815
R1326 AVSS.n1753 AVSS.n17 218.815
R1327 AVSS.n1753 AVSS.n26 218.815
R1328 AVSS.n1753 AVSS.n31 218.815
R1329 AVSS.n1753 AVSS.n36 218.815
R1330 AVSS.n1753 AVSS.n16 200.267
R1331 AVSS.n39 AVSS.n16 184.47
R1332 AVSS.n19 AVSS.n16 184.47
R1333 AVSS.n407 AVSS.n406 147.374
R1334 AVSS.n634 AVSS.n403 147.374
R1335 AVSS.n632 AVSS.n631 147.374
R1336 AVSS.n416 AVSS.n415 147.374
R1337 AVSS.n622 AVSS.n621 147.374
R1338 AVSS.n609 AVSS.n423 147.374
R1339 AVSS.n607 AVSS.n606 147.374
R1340 AVSS.n599 AVSS.n432 147.374
R1341 AVSS.n597 AVSS.n596 147.374
R1342 AVSS.n589 AVSS.n440 147.374
R1343 AVSS.n587 AVSS.n586 147.374
R1344 AVSS.n458 AVSS.n455 147.374
R1345 AVSS.n576 AVSS.n460 147.374
R1346 AVSS.n574 AVSS.n573 147.374
R1347 AVSS.n566 AVSS.n468 147.374
R1348 AVSS.n564 AVSS.n563 147.374
R1349 AVSS.n555 AVSS.n483 147.374
R1350 AVSS.n553 AVSS.n552 147.374
R1351 AVSS.n545 AVSS.n491 147.374
R1352 AVSS.n543 AVSS.n542 147.374
R1353 AVSS.n534 AVSS.n499 147.374
R1354 AVSS.n532 AVSS.n531 147.374
R1355 AVSS.n519 AVSS.n507 147.374
R1356 AVSS.n517 AVSS.n516 147.374
R1357 AVSS.n1683 AVSS.n1682 147.374
R1358 AVSS.n1406 AVSS.n1405 147.374
R1359 AVSS.n1409 AVSS.n1408 147.374
R1360 AVSS.n1418 AVSS.n1417 147.374
R1361 AVSS.n1421 AVSS.n1420 147.374
R1362 AVSS.n1434 AVSS.n1433 147.374
R1363 AVSS.n1437 AVSS.n1436 147.374
R1364 AVSS.n1447 AVSS.n1446 147.374
R1365 AVSS.n1450 AVSS.n1449 147.374
R1366 AVSS.n1461 AVSS.n1460 147.374
R1367 AVSS.n1464 AVSS.n1463 147.374
R1368 AVSS.n1367 AVSS.n1364 147.374
R1369 AVSS.n1477 AVSS.n1476 147.374
R1370 AVSS.n1480 AVSS.n1479 147.374
R1371 AVSS.n1496 AVSS.n1495 147.374
R1372 AVSS.n1499 AVSS.n1498 147.374
R1373 AVSS.n1510 AVSS.n1509 147.374
R1374 AVSS.n1513 AVSS.n1512 147.374
R1375 AVSS.n1521 AVSS.n1520 147.374
R1376 AVSS.n1339 AVSS.n1338 147.374
R1377 AVSS.n1533 AVSS.n1532 147.374
R1378 AVSS.n1536 AVSS.n1535 147.374
R1379 AVSS.n1548 AVSS.n1547 147.374
R1380 AVSS.n1551 AVSS.n1550 147.374
R1381 AVSS.n1669 AVSS.n1668 147.374
R1382 AVSS.n1672 AVSS.n1671 147.374
R1383 AVSS.n1684 AVSS.n1683 147.374
R1384 AVSS.n1407 AVSS.n1406 147.374
R1385 AVSS.n1408 AVSS.n1390 147.374
R1386 AVSS.n1419 AVSS.n1418 147.374
R1387 AVSS.n1420 AVSS.n1380 147.374
R1388 AVSS.n1435 AVSS.n1434 147.374
R1389 AVSS.n1436 AVSS.n1375 147.374
R1390 AVSS.n1448 AVSS.n1447 147.374
R1391 AVSS.n1449 AVSS.n1370 147.374
R1392 AVSS.n1462 AVSS.n1461 147.374
R1393 AVSS.n1465 AVSS.n1464 147.374
R1394 AVSS.n1364 AVSS.n1355 147.374
R1395 AVSS.n1478 AVSS.n1477 147.374
R1396 AVSS.n1479 AVSS.n1350 147.374
R1397 AVSS.n1497 AVSS.n1496 147.374
R1398 AVSS.n1498 AVSS.n1345 147.374
R1399 AVSS.n1511 AVSS.n1510 147.374
R1400 AVSS.n1512 AVSS.n1340 147.374
R1401 AVSS.n1522 AVSS.n1521 147.374
R1402 AVSS.n1338 AVSS.n1334 147.374
R1403 AVSS.n1534 AVSS.n1533 147.374
R1404 AVSS.n1535 AVSS.n1324 147.374
R1405 AVSS.n1549 AVSS.n1548 147.374
R1406 AVSS.n1550 AVSS.n1319 147.374
R1407 AVSS.n1670 AVSS.n1669 147.374
R1408 AVSS.n1671 AVSS.n1311 147.374
R1409 AVSS.n518 AVSS.n517 147.374
R1410 AVSS.n507 AVSS.n500 147.374
R1411 AVSS.n533 AVSS.n532 147.374
R1412 AVSS.n499 AVSS.n493 147.374
R1413 AVSS.n544 AVSS.n543 147.374
R1414 AVSS.n491 AVSS.n485 147.374
R1415 AVSS.n554 AVSS.n553 147.374
R1416 AVSS.n483 AVSS.n470 147.374
R1417 AVSS.n565 AVSS.n564 147.374
R1418 AVSS.n468 AVSS.n462 147.374
R1419 AVSS.n575 AVSS.n574 147.374
R1420 AVSS.n460 AVSS.n459 147.374
R1421 AVSS.n455 AVSS.n442 147.374
R1422 AVSS.n588 AVSS.n587 147.374
R1423 AVSS.n440 AVSS.n434 147.374
R1424 AVSS.n598 AVSS.n597 147.374
R1425 AVSS.n432 AVSS.n425 147.374
R1426 AVSS.n608 AVSS.n607 147.374
R1427 AVSS.n423 AVSS.n417 147.374
R1428 AVSS.n623 AVSS.n622 147.374
R1429 AVSS.n415 AVSS.n409 147.374
R1430 AVSS.n633 AVSS.n632 147.374
R1431 AVSS.n405 AVSS.n403 147.374
R1432 AVSS.n407 AVSS.n393 147.374
R1433 AVSS.n1752 AVSS.n1751 147.374
R1434 AVSS.n20 AVSS.n17 147.374
R1435 AVSS.n26 AVSS.n25 147.374
R1436 AVSS.n31 AVSS.n30 147.374
R1437 AVSS.n36 AVSS.n35 147.374
R1438 AVSS.n906 AVSS.n905 147.374
R1439 AVSS.n888 AVSS.n292 147.374
R1440 AVSS.n892 AVSS.n891 147.374
R1441 AVSS.n895 AVSS.n894 147.374
R1442 AVSS.n886 AVSS.n884 147.374
R1443 AVSS.n881 AVSS.n879 147.374
R1444 AVSS.n876 AVSS.n874 147.374
R1445 AVSS.n874 AVSS.n873 147.374
R1446 AVSS.n879 AVSS.n878 147.374
R1447 AVSS.n884 AVSS.n883 147.374
R1448 AVSS.n896 AVSS.n895 147.374
R1449 AVSS.n893 AVSS.n892 147.374
R1450 AVSS.n889 AVSS.n888 147.374
R1451 AVSS.n905 AVSS.n904 147.374
R1452 AVSS.n1752 AVSS.n41 147.374
R1453 AVSS.n23 AVSS.n17 147.374
R1454 AVSS.n28 AVSS.n26 147.374
R1455 AVSS.n33 AVSS.n31 147.374
R1456 AVSS.n36 AVSS.n13 147.374
R1457 AVSS.n387 AVSS.n384 135.992
R1458 AVSS.n646 AVSS.n645 132.142
R1459 AVSS.n1691 AVSS.n1690 117.46
R1460 AVSS.n1218 AVSS.n43 117.46
R1461 AVSS.n369 AVSS.t111 114.441
R1462 AVSS.n428 AVSS.t17 114.441
R1463 AVSS.n445 AVSS.t177 114.441
R1464 AVSS.n559 AVSS.t73 114.441
R1465 AVSS.n538 AVSS.t137 114.441
R1466 AVSS.n1298 AVSS.t47 114.441
R1467 AVSS.n1429 AVSS.t97 114.441
R1468 AVSS.n1456 AVSS.t92 114.441
R1469 AVSS.n1504 AVSS.t140 114.441
R1470 AVSS.n1526 AVSS.t121 114.441
R1471 AVSS.n369 AVSS.t117 114.439
R1472 AVSS.n428 AVSS.t23 114.439
R1473 AVSS.n445 AVSS.t14 114.439
R1474 AVSS.n559 AVSS.t79 114.439
R1475 AVSS.n538 AVSS.t21 114.439
R1476 AVSS.n1298 AVSS.t58 114.439
R1477 AVSS.n1429 AVSS.t103 114.439
R1478 AVSS.n1456 AVSS.t95 114.439
R1479 AVSS.n1504 AVSS.t143 114.439
R1480 AVSS.n1526 AVSS.t168 114.439
R1481 AVSS.n1567 AVSS.t64 114.439
R1482 AVSS.n1677 AVSS.n1313 114.072
R1483 AVSS.n910 AVSS.n908 106.541
R1484 AVSS.n1755 AVSS.n12 106.541
R1485 AVSS.n408 AVSS.n392 103.495
R1486 AVSS.n1113 AVSS.t84 103.459
R1487 AVSS.n1111 AVSS.t128 103.459
R1488 AVSS.n1663 AVSS.t55 103.459
R1489 AVSS.n1613 AVSS.t43 103.459
R1490 AVSS.n1599 AVSS.t105 103.459
R1491 AVSS.n1222 AVSS.t124 103.459
R1492 AVSS.n99 AVSS.t81 103.459
R1493 AVSS.n1051 AVSS.t39 103.459
R1494 AVSS.n209 AVSS.t160 103.459
R1495 AVSS.n974 AVSS.t51 103.459
R1496 AVSS.n917 AVSS.t61 103.459
R1497 AVSS.n724 AVSS.t25 103.459
R1498 AVSS.n295 AVSS.t29 103.459
R1499 AVSS.n667 AVSS.t114 103.459
R1500 AVSS.n385 AVSS.t119 103.459
R1501 AVSS.n94 AVSS.t100 103.459
R1502 AVSS.n1146 AVSS.t134 103.459
R1503 AVSS.n163 AVSS.t66 103.459
R1504 AVSS.n206 AVSS.t71 103.459
R1505 AVSS.n1010 AVSS.t163 103.459
R1506 AVSS.n284 AVSS.t32 103.459
R1507 AVSS.n867 AVSS.t174 103.459
R1508 AVSS.n795 AVSS.t76 103.459
R1509 AVSS.n1132 AVSS.t11 103.459
R1510 AVSS.n828 AVSS.t88 103.459
R1511 AVSS.n839 AVSS.t90 103.459
R1512 AVSS.n846 AVSS.t36 103.459
R1513 AVSS.n1715 AVSS.t149 103.459
R1514 AVSS.n1261 AVSS.t68 103.459
R1515 AVSS.n1203 AVSS.t170 103.459
R1516 AVSS.n79 AVSS.t108 103.459
R1517 AVSS.n1081 AVSS.t145 103.459
R1518 AVSS.n188 AVSS.t153 103.459
R1519 AVSS.n961 AVSS.t156 103.459
R1520 AVSS.n937 AVSS.t165 103.459
R1521 AVSS.n321 AVSS.t7 103.459
R1522 AVSS.n707 AVSS.t131 103.459
R1523 AVSS.n872 AVSS.n871 101.272
R1524 AVSS.n1680 AVSS.n1306 93.855
R1525 AVSS.n224 AVSS.t195 87.245
R1526 AVSS.n225 AVSS.t190 87.245
R1527 AVSS.n226 AVSS.t183 87.245
R1528 AVSS.n227 AVSS.t187 87.245
R1529 AVSS.n1586 AVSS.t193 87.2444
R1530 AVSS.n1585 AVSS.t196 87.2444
R1531 AVSS.n1584 AVSS.t181 87.2444
R1532 AVSS.n1583 AVSS.t205 87.2444
R1533 AVSS.n1586 AVSS.t206 87.2437
R1534 AVSS.n1585 AVSS.t186 87.2437
R1535 AVSS.n1584 AVSS.t200 87.2437
R1536 AVSS.n1583 AVSS.t201 87.2437
R1537 AVSS.n224 AVSS.t203 87.2431
R1538 AVSS.n225 AVSS.t189 87.2431
R1539 AVSS.n226 AVSS.t197 87.2431
R1540 AVSS.n227 AVSS.t198 87.2431
R1541 AVSS.n503 AVSS.t199 87.2137
R1542 AVSS.n474 AVSS.t192 87.2137
R1543 AVSS.n448 AVSS.t204 87.2137
R1544 AVSS.n617 AVSS.t202 87.2137
R1545 AVSS.n1105 AVSS.t6 87.1994
R1546 AVSS.n0 AVSS.t87 87.1387
R1547 AVSS.n1106 AVSS.t86 87.1387
R1548 AVSS.n1314 AVSS.t57 87.1387
R1549 AVSS.t65 AVSS.n1642 87.1387
R1550 AVSS.n1623 AVSS.t46 87.1387
R1551 AVSS.t107 AVSS.n1609 87.1387
R1552 AVSS.n45 AVSS.t127 87.1387
R1553 AVSS.n1178 AVSS.t83 87.1387
R1554 AVSS.n1063 AVSS.t42 87.1387
R1555 AVSS.n1014 AVSS.t162 87.1387
R1556 AVSS.n976 AVSS.t54 87.1387
R1557 AVSS.t63 AVSS.n925 87.1387
R1558 AVSS.n731 AVSS.t28 87.1387
R1559 AVSS.t31 AVSS.n718 87.1387
R1560 AVSS.n670 AVSS.t116 87.1387
R1561 AVSS.t120 AVSS.n655 87.1387
R1562 AVSS.n62 AVSS.t102 87.1387
R1563 AVSS.n1186 AVSS.t101 87.1387
R1564 AVSS.n1155 AVSS.t136 87.1387
R1565 AVSS.n247 AVSS.t164 87.1387
R1566 AVSS.n255 AVSS.t35 87.1387
R1567 AVSS.n919 AVSS.t34 87.1387
R1568 AVSS.n797 AVSS.t176 87.1387
R1569 AVSS.n787 AVSS.t175 87.1387
R1570 AVSS.n1100 AVSS.t13 87.1387
R1571 AVSS.t38 AVSS.n818 87.1387
R1572 AVSS.n1282 AVSS.t152 87.1387
R1573 AVSS.t70 AVSS.n1248 87.1387
R1574 AVSS.n1235 AVSS.t173 87.1387
R1575 AVSS.t110 AVSS.n1197 87.1387
R1576 AVSS.n1086 AVSS.t148 87.1387
R1577 AVSS.t155 AVSS.n1032 87.1387
R1578 AVSS.n957 AVSS.t159 87.1387
R1579 AVSS.t167 AVSS.n952 87.1387
R1580 AVSS.n760 AVSS.t10 87.1387
R1581 AVSS.n704 AVSS.t133 87.1387
R1582 AVSS.n0 AVSS.t130 87.1377
R1583 AVSS.n1106 AVSS.t129 87.1377
R1584 AVSS.n797 AVSS.t78 87.1377
R1585 AVSS.n787 AVSS.t77 87.1377
R1586 AVSS.n639 AVSS.t113 76.1469
R1587 AVSS.n398 AVSS.t118 76.1469
R1588 AVSS.n615 AVSS.t20 76.1469
R1589 AVSS.n614 AVSS.t24 76.1469
R1590 AVSS.n581 AVSS.t179 76.1469
R1591 AVSS.n450 AVSS.t16 76.1469
R1592 AVSS.n478 AVSS.t75 76.1469
R1593 AVSS.n477 AVSS.t80 76.1469
R1594 AVSS.n526 AVSS.t139 76.1469
R1595 AVSS.n524 AVSS.t22 76.1469
R1596 AVSS.n1399 AVSS.t50 76.1469
R1597 AVSS.n1398 AVSS.t60 76.1469
R1598 AVSS.n1426 AVSS.t99 76.1469
R1599 AVSS.n1385 AVSS.t104 76.1469
R1600 AVSS.n1470 AVSS.t94 76.1469
R1601 AVSS.n1360 AVSS.t96 76.1469
R1602 AVSS.n1490 AVSS.t142 76.1469
R1603 AVSS.n1489 AVSS.t144 76.1469
R1604 AVSS.n1541 AVSS.t123 76.1469
R1605 AVSS.n1329 AVSS.t169 76.1469
R1606 AVSS.n1644 AVSS.n1643 69.7387
R1607 AVSS.n1611 AVSS.n1610 69.7387
R1608 AVSS.n1177 AVSS.n65 69.7387
R1609 AVSS.n1013 AVSS.n168 69.7387
R1610 AVSS.n927 AVSS.n926 69.7387
R1611 AVSS.n720 AVSS.n719 69.7387
R1612 AVSS.n657 AVSS.n656 69.7387
R1613 AVSS.n1062 AVSS.n1060 69.7387
R1614 AVSS.n1059 AVSS.n1058 69.7387
R1615 AVSS.n240 AVSS.n200 69.7387
R1616 AVSS.n820 AVSS.n135 69.7387
R1617 AVSS.n822 AVSS.n821 69.7387
R1618 AVSS.n819 AVSS.n807 69.7387
R1619 AVSS.n1265 AVSS.n1264 69.7387
R1620 AVSS.n1199 AVSS.n1198 69.7387
R1621 AVSS.n1034 AVSS.n1033 69.7387
R1622 AVSS.n954 AVSS.n953 69.7387
R1623 AVSS.n772 AVSS.n308 69.7387
R1624 AVSS.n397 AVSS.n395 58.7469
R1625 AVSS.n613 AVSS.n420 58.7469
R1626 AVSS.n449 AVSS.n447 58.7469
R1627 AVSS.n476 AVSS.n475 58.7469
R1628 AVSS.n523 AVSS.n504 58.7469
R1629 AVSS.n1397 AVSS.n1396 58.7469
R1630 AVSS.n1384 AVSS.n1383 58.7469
R1631 AVSS.n1359 AVSS.n1358 58.7469
R1632 AVSS.n1488 AVSS.n1487 58.7469
R1633 AVSS.n1328 AVSS.n1327 58.7469
R1634 AVSS.n650 AVSS.n392 34.4984
R1635 AVSS.n682 AVSS.n374 34.4984
R1636 AVSS.n682 AVSS.n681 34.4984
R1637 AVSS.n680 AVSS.n675 34.4984
R1638 AVSS.n675 AVSS.n355 34.4984
R1639 AVSS.n690 AVSS.n355 34.4984
R1640 AVSS.n690 AVSS.n356 34.4984
R1641 AVSS.n356 AVSS.n348 34.4984
R1642 AVSS.n700 AVSS.n348 34.4984
R1643 AVSS.n700 AVSS.n340 34.4984
R1644 AVSS.n713 AVSS.n340 34.4984
R1645 AVSS.n777 AVSS.n301 34.4984
R1646 AVSS.n777 AVSS.n302 34.4984
R1647 AVSS.n767 AVSS.n302 34.4984
R1648 AVSS.n766 AVSS.n765 34.4984
R1649 AVSS.n765 AVSS.n315 34.4984
R1650 AVSS.n755 AVSS.n315 34.4984
R1651 AVSS.n755 AVSS.n754 34.4984
R1652 AVSS.n754 AVSS.n753 34.4984
R1653 AVSS.n753 AVSS.n746 34.4984
R1654 AVSS.n947 AVSS.n946 34.4984
R1655 AVSS.n1740 AVSS.n37 34.4984
R1656 AVSS.n1740 AVSS.n51 34.4984
R1657 AVSS.n1734 AVSS.n51 34.4984
R1658 AVSS.n1734 AVSS.n1733 34.4984
R1659 AVSS.n1733 AVSS.n1732 34.4984
R1660 AVSS.n1732 AVSS.n1243 34.4984
R1661 AVSS.n1722 AVSS.n1721 34.4984
R1662 AVSS.n1721 AVSS.n1255 34.4984
R1663 AVSS.n1709 AVSS.n1273 34.4984
R1664 AVSS.n1709 AVSS.n1708 34.4984
R1665 AVSS.n1708 AVSS.n1707 34.4984
R1666 AVSS.n1707 AVSS.n1277 34.4984
R1667 AVSS.n1698 AVSS.n1277 34.4984
R1668 AVSS.n1698 AVSS.n1697 34.4984
R1669 AVSS.n1697 AVSS.n1696 34.4984
R1670 AVSS.n1696 AVSS.n1290 34.4984
R1671 AVSS.n1649 AVSS.n1561 34.4984
R1672 AVSS.n1649 AVSS.n1558 34.4984
R1673 AVSS.n1655 AVSS.n1558 34.4984
R1674 AVSS.n1680 AVSS.n1309 34.4984
R1675 AVSS.n510 AVSS.n384 34.3446
R1676 AVSS.n681 AVSS.t18 33.4837
R1677 AVSS.t69 AVSS.n1722 33.4837
R1678 AVSS.n788 AVSS.n293 33.1299
R1679 AVSS.n38 AVSS.n7 33.1299
R1680 AVSS.t180 AVSS.n1243 31.4544
R1681 AVSS.n746 AVSS.n272 30.9471
R1682 AVSS.n933 AVSS.n276 30.9471
R1683 AVSS.n967 AVSS.n260 30.9471
R1684 AVSS.n982 AVSS.n981 30.9471
R1685 AVSS.n993 AVSS.n231 30.9471
R1686 AVSS.n992 AVSS.n234 30.9471
R1687 AVSS.n1005 AVSS.n218 30.9471
R1688 AVSS.n1026 AVSS.n192 30.9471
R1689 AVSS.n1025 AVSS.n195 30.9471
R1690 AVSS.n180 AVSS.n172 30.9471
R1691 AVSS.n1049 AVSS.n1048 30.9471
R1692 AVSS.n1074 AVSS.n148 30.9471
R1693 AVSS.n1091 AVSS.n138 30.9471
R1694 AVSS.n1092 AVSS.n130 30.9471
R1695 AVSS.n1140 AVSS.n1139 30.9471
R1696 AVSS.n1161 AVSS.n116 30.9471
R1697 AVSS.n1172 AVSS.n106 30.9471
R1698 AVSS.n108 AVSS.n107 30.9471
R1699 AVSS.n1192 AVSS.n84 30.9471
R1700 AVSS.n1209 AVSS.n68 30.9471
R1701 AVSS.n1228 AVSS.n59 30.9471
R1702 AVSS.t15 AVSS.n374 28.4105
R1703 AVSS.t157 AVSS.n250 28.4105
R1704 AVSS.t37 AVSS.n219 28.4105
R1705 AVSS.n1753 AVSS.n15 28.4105
R1706 AVSS.t85 AVSS.n69 27.9032
R1707 AVSS.n514 AVSS.n510 27.1064
R1708 AVSS.n702 AVSS.n345 25.6005
R1709 AVSS.n702 AVSS.n346 25.6005
R1710 AVSS.n941 AVSS.n263 25.6005
R1711 AVSS.n965 AVSS.n263 25.6005
R1712 AVSS.n184 AVSS.n146 25.6005
R1713 AVSS.n1076 AVSS.n146 25.6005
R1714 AVSS.n1738 AVSS.n1737 25.6005
R1715 AVSS.n1737 AVSS.n1736 25.6005
R1716 AVSS.n1297 AVSS.n1294 25.6005
R1717 AVSS.n1560 AVSS.n1297 25.6005
R1718 AVSS.n630 AVSS.n629 25.6005
R1719 AVSS.n457 AVSS.n453 25.6005
R1720 AVSS.n535 AVSS.n498 25.6005
R1721 AVSS.n698 AVSS.n697 25.6005
R1722 AVSS.n698 AVSS.n337 25.6005
R1723 AVSS.n912 AVSS.n258 25.6005
R1724 AVSS.n969 AVSS.n258 25.6005
R1725 AVSS.n1056 AVSS.n170 25.6005
R1726 AVSS.n1056 AVSS.n1055 25.6005
R1727 AVSS.n1588 AVSS.n50 25.6005
R1728 AVSS.n1588 AVSS.n1579 25.6005
R1729 AVSS.n1637 AVSS.n1563 25.6005
R1730 AVSS.n1647 AVSS.n1563 25.6005
R1731 AVSS.n1410 AVSS.n1391 25.6005
R1732 AVSS.n1366 AVSS.n1365 25.6005
R1733 AVSS.n1531 AVSS.n1331 25.6005
R1734 AVSS.n887 AVSS.n792 25.6005
R1735 AVSS.n979 AVSS.n253 25.6005
R1736 AVSS.n124 AVSS.n123 25.6005
R1737 AVSS.n22 AVSS.n21 25.6005
R1738 AVSS.n863 AVSS.n860 25.6005
R1739 AVSS.n1129 AVSS.n1101 25.6005
R1740 AVSS.n713 AVSS.t191 25.3666
R1741 AVSS.t171 AVSS.n15 25.3666
R1742 AVSS.t48 AVSS.n1309 25.3666
R1743 AVSS.n410 AVSS.n404 25.224
R1744 AVSS.n456 AVSS.n444 25.224
R1745 AVSS.n536 AVSS.n495 25.224
R1746 AVSS.n1411 AVSS.n1393 25.224
R1747 AVSS.n1466 AVSS.n1363 25.224
R1748 AVSS.n1530 AVSS.n1529 25.224
R1749 AVSS.n890 AVSS.n786 25.224
R1750 AVSS.n978 AVSS.n254 25.224
R1751 AVSS.n121 AVSS.n120 25.224
R1752 AVSS.n18 AVSS.n5 25.224
R1753 AVSS.n859 AVSS.n801 25.224
R1754 AVSS.n1125 AVSS.n1102 25.224
R1755 AVSS.n812 AVSS.t182 24.8593
R1756 AVSS.n628 AVSS.n411 24.4711
R1757 AVSS.n578 AVSS.n577 24.4711
R1758 AVSS.n530 AVSS.n501 24.4711
R1759 AVSS.n1416 AVSS.n1414 24.4711
R1760 AVSS.n1475 AVSS.n1356 24.4711
R1761 AVSS.n1538 AVSS.n1537 24.4711
R1762 AVSS.n898 AVSS.n897 24.4711
R1763 AVSS.n283 AVSS.n257 24.4711
R1764 AVSS.n1159 AVSS.n1158 24.4711
R1765 AVSS.n24 AVSS.n8 24.4711
R1766 AVSS.n864 AVSS.n799 24.4711
R1767 AVSS.n1130 AVSS.n134 24.4711
R1768 AVSS.t194 AVSS.n1255 24.3519
R1769 AVSS.n363 AVSS.n360 24.0946
R1770 AVSS.n711 AVSS.n342 24.0946
R1771 AVSS.n943 AVSS.n942 24.0946
R1772 AVSS.n964 AVSS.n264 24.0946
R1773 AVSS.n1037 AVSS.n1036 24.0946
R1774 AVSS.n1078 AVSS.n1077 24.0946
R1775 AVSS.n1232 AVSS.n54 24.0946
R1776 AVSS.n1245 AVSS.n1238 24.0946
R1777 AVSS.n1694 AVSS.n1693 24.0946
R1778 AVSS.n1651 AVSS.n1299 24.0946
R1779 AVSS.n696 AVSS.n350 24.0946
R1780 AVSS.n716 AVSS.n715 24.0946
R1781 AVSS.n914 AVSS.n913 24.0946
R1782 AVSS.n971 AVSS.n970 24.0946
R1783 AVSS.n1042 AVSS.n1041 24.0946
R1784 AVSS.n1054 AVSS.n159 24.0946
R1785 AVSS.n1743 AVSS.n47 24.0946
R1786 AVSS.n1593 AVSS.n1592 24.0946
R1787 AVSS.n1639 AVSS.n1638 24.0946
R1788 AVSS.n1646 AVSS.n1564 24.0946
R1789 AVSS.n635 AVSS.n402 23.7181
R1790 AVSS.n585 AVSS.n584 23.7181
R1791 AVSS.n541 AVSS.n540 23.7181
R1792 AVSS.n1404 AVSS.n1403 23.7181
R1793 AVSS.n1467 AVSS.n1362 23.7181
R1794 AVSS.n1528 AVSS.n1335 23.7181
R1795 AVSS.n990 AVSS.n237 23.7181
R1796 AVSS.n1189 AVSS.n91 23.7181
R1797 AVSS.n856 AVSS.n855 23.7181
R1798 AVSS.n1124 AVSS.n1103 23.7181
R1799 AVSS.n625 AVSS.n624 22.9652
R1800 AVSS.n461 AVSS.n454 22.9652
R1801 AVSS.n529 AVSS.n502 22.9652
R1802 AVSS.n1415 AVSS.n1387 22.9652
R1803 AVSS.n1474 AVSS.n1354 22.9652
R1804 AVSS.n1333 AVSS.n1332 22.9652
R1805 AVSS.n885 AVSS.n783 22.9652
R1806 AVSS.n930 AVSS.n929 22.9652
R1807 AVSS.n1143 AVSS.n119 22.9652
R1808 AVSS.n27 AVSS.n3 22.9652
R1809 AVSS.n798 AVSS.n794 22.9652
R1810 AVSS.n1136 AVSS.n1135 22.9652
R1811 AVSS.n688 AVSS.n687 22.5887
R1812 AVSS.n710 AVSS.n343 22.5887
R1813 AVSS.n940 AVSS.n935 22.5887
R1814 AVSS.n959 AVSS.n958 22.5887
R1815 AVSS.n1029 AVSS.n183 22.5887
R1816 AVSS.n1089 AVSS.n142 22.5887
R1817 AVSS.n1233 AVSS.n1231 22.5887
R1818 AVSS.n1730 AVSS.n1246 22.5887
R1819 AVSS.n1293 AVSS.n1292 22.5887
R1820 AVSS.n1653 AVSS.n1296 22.5887
R1821 AVSS.n693 AVSS.n692 22.5887
R1822 AVSS.n338 AVSS.n297 22.5887
R1823 AVSS.n915 AVSS.n289 22.5887
R1824 AVSS.n984 AVSS.n248 22.5887
R1825 AVSS.n1018 AVSS.n178 22.5887
R1826 AVSS.n1067 AVSS.n1066 22.5887
R1827 AVSS.n1744 AVSS.n46 22.5887
R1828 AVSS.n1595 AVSS.n1594 22.5887
R1829 AVSS.n1640 AVSS.n1635 22.5887
R1830 AVSS.n1657 AVSS.n1556 22.5887
R1831 AVSS.n901 AVSS.n900 22.5887
R1832 AVSS.n1746 AVSS.n4 22.5887
R1833 AVSS.n636 AVSS.n401 22.2123
R1834 AVSS.n443 AVSS.n441 22.2123
R1835 AVSS.n494 AVSS.n492 22.2123
R1836 AVSS.n1402 AVSS.n1394 22.2123
R1837 AVSS.n1369 AVSS.n1368 22.2123
R1838 AVSS.n1524 AVSS.n1523 22.2123
R1839 AVSS.n989 AVSS.n238 22.2123
R1840 AVSS.n1188 AVSS.n92 22.2123
R1841 AVSS.n854 AVSS.n853 22.2123
R1842 AVSS.n1121 AVSS.n1120 22.2123
R1843 AVSS.n640 AVSS.n639 21.9824
R1844 AVSS.n640 AVSS.n395 21.9824
R1845 AVSS.n640 AVSS.n398 21.9824
R1846 AVSS.n615 AVSS.n419 21.9824
R1847 AVSS.n420 AVSS.n419 21.9824
R1848 AVSS.n614 AVSS.n419 21.9824
R1849 AVSS.n582 AVSS.n581 21.9824
R1850 AVSS.n582 AVSS.n447 21.9824
R1851 AVSS.n582 AVSS.n450 21.9824
R1852 AVSS.n478 AVSS.n466 21.9824
R1853 AVSS.n475 AVSS.n466 21.9824
R1854 AVSS.n477 AVSS.n466 21.9824
R1855 AVSS.n526 AVSS.n525 21.9824
R1856 AVSS.n525 AVSS.n504 21.9824
R1857 AVSS.n525 AVSS.n524 21.9824
R1858 AVSS.n1399 AVSS.n1303 21.9824
R1859 AVSS.n1396 AVSS.n1303 21.9824
R1860 AVSS.n1398 AVSS.n1303 21.9824
R1861 AVSS.n1426 AVSS.n1425 21.9824
R1862 AVSS.n1425 AVSS.n1383 21.9824
R1863 AVSS.n1425 AVSS.n1385 21.9824
R1864 AVSS.n1470 AVSS.n1469 21.9824
R1865 AVSS.n1469 AVSS.n1358 21.9824
R1866 AVSS.n1469 AVSS.n1360 21.9824
R1867 AVSS.n1490 AVSS.n1486 21.9824
R1868 AVSS.n1487 AVSS.n1486 21.9824
R1869 AVSS.n1489 AVSS.n1486 21.9824
R1870 AVSS.n1541 AVSS.n1540 21.9824
R1871 AVSS.n1540 AVSS.n1327 21.9824
R1872 AVSS.n1540 AVSS.n1329 21.9824
R1873 AVSS.n639 AVSS.n638 21.982
R1874 AVSS.n638 AVSS.n395 21.982
R1875 AVSS.n638 AVSS.n398 21.982
R1876 AVSS.n616 AVSS.n615 21.982
R1877 AVSS.n616 AVSS.n420 21.982
R1878 AVSS.n616 AVSS.n614 21.982
R1879 AVSS.n581 AVSS.n580 21.982
R1880 AVSS.n580 AVSS.n447 21.982
R1881 AVSS.n580 AVSS.n450 21.982
R1882 AVSS.n479 AVSS.n478 21.982
R1883 AVSS.n479 AVSS.n475 21.982
R1884 AVSS.n479 AVSS.n477 21.982
R1885 AVSS.n527 AVSS.n526 21.982
R1886 AVSS.n527 AVSS.n504 21.982
R1887 AVSS.n527 AVSS.n524 21.982
R1888 AVSS.n1400 AVSS.n1399 21.982
R1889 AVSS.n1400 AVSS.n1396 21.982
R1890 AVSS.n1400 AVSS.n1398 21.982
R1891 AVSS.n1427 AVSS.n1426 21.982
R1892 AVSS.n1427 AVSS.n1383 21.982
R1893 AVSS.n1427 AVSS.n1385 21.982
R1894 AVSS.n1471 AVSS.n1470 21.982
R1895 AVSS.n1471 AVSS.n1358 21.982
R1896 AVSS.n1471 AVSS.n1360 21.982
R1897 AVSS.n1491 AVSS.n1490 21.982
R1898 AVSS.n1491 AVSS.n1487 21.982
R1899 AVSS.n1491 AVSS.n1489 21.982
R1900 AVSS.n1542 AVSS.n1541 21.982
R1901 AVSS.n1542 AVSS.n1327 21.982
R1902 AVSS.n1542 AVSS.n1329 21.982
R1903 AVSS.n1113 AVSS.n1110 21.9607
R1904 AVSS.n1114 AVSS.n1113 21.9607
R1905 AVSS.n1111 AVSS.n1110 21.9607
R1906 AVSS.n1114 AVSS.n1111 21.9607
R1907 AVSS.n1664 AVSS.n1663 21.9607
R1908 AVSS.n1663 AVSS.n1662 21.9607
R1909 AVSS.n1614 AVSS.n1613 21.9607
R1910 AVSS.n1613 AVSS.n1573 21.9607
R1911 AVSS.n1599 AVSS.n1598 21.9607
R1912 AVSS.n1600 AVSS.n1599 21.9607
R1913 AVSS.n1222 AVSS.n1221 21.9607
R1914 AVSS.n1223 AVSS.n1222 21.9607
R1915 AVSS.n99 AVSS.n93 21.9607
R1916 AVSS.n100 AVSS.n99 21.9607
R1917 AVSS.n1052 AVSS.n1051 21.9607
R1918 AVSS.n1051 AVSS.n156 21.9607
R1919 AVSS.n210 AVSS.n209 21.9607
R1920 AVSS.n209 AVSS.n208 21.9607
R1921 AVSS.n974 AVSS.n973 21.9607
R1922 AVSS.n975 AVSS.n974 21.9607
R1923 AVSS.n917 AVSS.n290 21.9607
R1924 AVSS.n918 AVSS.n917 21.9607
R1925 AVSS.n725 AVSS.n724 21.9607
R1926 AVSS.n724 AVSS.n332 21.9607
R1927 AVSS.n295 AVSS.n294 21.9607
R1928 AVSS.n296 AVSS.n295 21.9607
R1929 AVSS.n667 AVSS.n666 21.9607
R1930 AVSS.n668 AVSS.n667 21.9607
R1931 AVSS.n386 AVSS.n385 21.9607
R1932 AVSS.n385 AVSS.n383 21.9607
R1933 AVSS.n95 AVSS.n94 21.9607
R1934 AVSS.n94 AVSS.n63 21.9607
R1935 AVSS.n1147 AVSS.n1146 21.9607
R1936 AVSS.n1146 AVSS.n125 21.9607
R1937 AVSS.n163 AVSS.n155 21.9607
R1938 AVSS.n164 AVSS.n163 21.9607
R1939 AVSS.n206 AVSS.n201 21.9607
R1940 AVSS.n207 AVSS.n206 21.9607
R1941 AVSS.n1010 AVSS.n1009 21.9607
R1942 AVSS.n1011 AVSS.n1010 21.9607
R1943 AVSS.n285 AVSS.n284 21.9607
R1944 AVSS.n284 AVSS.n256 21.9607
R1945 AVSS.n868 AVSS.n867 21.9607
R1946 AVSS.n867 AVSS.n866 21.9607
R1947 AVSS.n868 AVSS.n795 21.9607
R1948 AVSS.n866 AVSS.n795 21.9607
R1949 AVSS.n1132 AVSS.n1099 21.9607
R1950 AVSS.n1133 AVSS.n1132 21.9607
R1951 AVSS.n829 AVSS.n828 21.9607
R1952 AVSS.n828 AVSS.n827 21.9607
R1953 AVSS.n840 AVSS.n839 21.9607
R1954 AVSS.n839 AVSS.n838 21.9607
R1955 AVSS.n846 AVSS.n806 21.9607
R1956 AVSS.n847 AVSS.n846 21.9607
R1957 AVSS.n1716 AVSS.n1715 21.9607
R1958 AVSS.n1715 AVSS.n1714 21.9607
R1959 AVSS.n1261 AVSS.n1249 21.9607
R1960 AVSS.n1262 AVSS.n1261 21.9607
R1961 AVSS.n1204 AVSS.n1203 21.9607
R1962 AVSS.n1203 AVSS.n1202 21.9607
R1963 AVSS.n79 AVSS.n76 21.9607
R1964 AVSS.n80 AVSS.n79 21.9607
R1965 AVSS.n1081 AVSS.n1080 21.9607
R1966 AVSS.n1082 AVSS.n1081 21.9607
R1967 AVSS.n189 AVSS.n188 21.9607
R1968 AVSS.n188 AVSS.n185 21.9607
R1969 AVSS.n961 AVSS.n956 21.9607
R1970 AVSS.n962 AVSS.n961 21.9607
R1971 AVSS.n937 AVSS.n936 21.9607
R1972 AVSS.n938 AVSS.n937 21.9607
R1973 AVSS.n321 AVSS.n309 21.9607
R1974 AVSS.n322 AVSS.n321 21.9607
R1975 AVSS.n708 AVSS.n707 21.9607
R1976 AVSS.n707 AVSS.n307 21.9607
R1977 AVSS.n620 AVSS.n414 21.4593
R1978 AVSS.n572 AVSS.n463 21.4593
R1979 AVSS.n521 AVSS.n520 21.4593
R1980 AVSS.n1423 AVSS.n1422 21.4593
R1981 AVSS.n1481 AVSS.n1353 21.4593
R1982 AVSS.n1546 AVSS.n1325 21.4593
R1983 AVSS.n882 AVSS.n791 21.4593
R1984 AVSS.n909 AVSS.n282 21.4593
R1985 AVSS.n1144 AVSS.n1142 21.4593
R1986 AVSS.n29 AVSS.n9 21.4593
R1987 AVSS.n871 AVSS.n870 21.4593
R1988 AVSS.n1095 AVSS.n133 21.4593
R1989 AVSS.t166 AVSS.n945 21.308
R1990 AVSS.n364 AVSS.n359 21.0829
R1991 AVSS.n775 AVSS.n305 21.0829
R1992 AVSS.n949 AVSS.n269 21.0829
R1993 AVSS.n995 AVSS.n229 21.0829
R1994 AVSS.n1030 AVSS.n1028 21.0829
R1995 AVSS.n1088 AVSS.n143 21.0829
R1996 AVSS.n58 AVSS.n56 21.0829
R1997 AVSS.n1729 AVSS.n1247 21.0829
R1998 AVSS.n1700 AVSS.n1285 21.0829
R1999 AVSS.n1307 AVSS.n1300 21.0829
R2000 AVSS.n379 AVSS.n352 21.0829
R2001 AVSS.n780 AVSS.n779 21.0829
R2002 AVSS.n922 AVSS.n921 21.0829
R2003 AVSS.n986 AVSS.n985 21.0829
R2004 AVSS.n1019 AVSS.n1017 21.0829
R2005 AVSS.n1065 AVSS.n162 21.0829
R2006 AVSS.n1226 AVSS.n1225 21.0829
R2007 AVSS.n1607 AVSS.n1606 21.0829
R2008 AVSS.n1634 AVSS.n1633 21.0829
R2009 AVSS.n1659 AVSS.n1658 21.0829
R2010 AVSS.n903 AVSS.n902 21.0829
R2011 AVSS.n1747 AVSS.n44 21.0829
R2012 AVSS.n400 AVSS.n394 20.7064
R2013 AVSS.n590 AVSS.n439 20.7064
R2014 AVSS.n546 AVSS.n490 20.7064
R2015 AVSS.n1685 AVSS.n1304 20.7064
R2016 AVSS.n1459 AVSS.n1458 20.7064
R2017 AVSS.n1519 AVSS.n1337 20.7064
R2018 AVSS.n245 AVSS.n244 20.7064
R2019 AVSS.n97 AVSS.n64 20.7064
R2020 AVSS.n850 AVSS.n803 20.7064
R2021 AVSS.n1117 AVSS.n1107 20.7064
R2022 AVSS.n619 AVSS.n418 19.9534
R2023 AVSS.n571 AVSS.n464 19.9534
R2024 AVSS.n508 AVSS.n506 19.9534
R2025 AVSS.n1389 AVSS.n1388 19.9534
R2026 AVSS.n1483 AVSS.n1482 19.9534
R2027 AVSS.n1545 AVSS.n1323 19.9534
R2028 AVSS.n880 AVSS.n784 19.9534
R2029 AVSS.n165 AVSS.n128 19.9534
R2030 AVSS.n32 AVSS.n2 19.9534
R2031 AVSS.n1096 AVSS.n1094 19.9534
R2032 AVSS.n676 AVSS.n365 19.577
R2033 AVSS.n774 AVSS.n306 19.577
R2034 AVSS.n950 AVSS.n268 19.577
R2035 AVSS.n997 AVSS.n996 19.577
R2036 AVSS.n223 AVSS.n190 19.577
R2037 AVSS.n1084 AVSS.n1083 19.577
R2038 AVSS.n1200 AVSS.n73 19.577
R2039 AVSS.n1726 AVSS.n1725 19.577
R2040 AVSS.n1701 AVSS.n1281 19.577
R2041 AVSS.n1301 AVSS.n1295 19.577
R2042 AVSS.n673 AVSS.n672 19.577
R2043 AVSS.n721 AVSS.n298 19.577
R2044 AVSS.n923 AVSS.n288 19.577
R2045 AVSS.n987 AVSS.n215 19.577
R2046 AVSS.n1016 AVSS.n211 19.577
R2047 AVSS.n160 AVSS.n126 19.577
R2048 AVSS.n1212 AVSS.n61 19.577
R2049 AVSS.n1604 AVSS.n1603 19.577
R2050 AVSS.n1632 AVSS.n1570 19.577
R2051 AVSS.n1678 AVSS.n1312 19.577
R2052 AVSS.n907 AVSS.n291 19.577
R2053 AVSS.n1750 AVSS.n1749 19.577
R2054 AVSS.n643 AVSS.n642 19.2005
R2055 AVSS.n591 AVSS.n436 19.2005
R2056 AVSS.n547 AVSS.n487 19.2005
R2057 AVSS.n1686 AVSS.n1302 19.2005
R2058 AVSS.n1452 AVSS.n1371 19.2005
R2059 AVSS.n1518 AVSS.n1341 19.2005
R2060 AVSS.n242 AVSS.n241 19.2005
R2061 AVSS.n1217 AVSS.n1216 19.2005
R2062 AVSS.n849 AVSS.n805 19.2005
R2063 AVSS.n1116 AVSS.n1108 19.2005
R2064 AVSS.n611 AVSS.n610 18.4476
R2065 AVSS.n568 AVSS.n567 18.4476
R2066 AVSS.n515 AVSS.n509 18.4476
R2067 AVSS.n1432 AVSS.n1381 18.4476
R2068 AVSS.n1494 AVSS.n1351 18.4476
R2069 AVSS.n1552 AVSS.n1322 18.4476
R2070 AVSS.n877 AVSS.n790 18.4476
R2071 AVSS.n166 AVSS.n154 18.4476
R2072 AVSS.n34 AVSS.n10 18.4476
R2073 AVSS.n823 AVSS.n136 18.4476
R2074 AVSS.n767 AVSS.t4 18.2641
R2075 AVSS.t109 AVSS.n87 18.2641
R2076 AVSS.n1561 AVSS.t59 18.2641
R2077 AVSS.n678 AVSS.n366 18.0711
R2078 AVSS.n770 AVSS.n769 18.0711
R2079 AVSS.n751 AVSS.n750 18.0711
R2080 AVSS.n1003 AVSS.n1002 18.0711
R2081 AVSS.n1164 AVSS.n112 18.0711
R2082 AVSS.n1207 AVSS.n1206 18.0711
R2083 AVSS.n1257 AVSS.n1250 18.0711
R2084 AVSS.n1705 AVSS.n1704 18.0711
R2085 AVSS.n661 AVSS.n378 18.0711
R2086 AVSS.n722 AVSS.n333 18.0711
R2087 AVSS.n743 AVSS.n742 18.0711
R2088 AVSS.n1007 AVSS.n213 18.0711
R2089 AVSS.n1151 AVSS.n1150 18.0711
R2090 AVSS.n1213 AVSS.n1211 18.0711
R2091 AVSS.n1602 AVSS.n1597 18.0711
R2092 AVSS.n1629 AVSS.n1628 18.0711
R2093 AVSS.n1073 AVSS.t2 17.7568
R2094 AVSS.n595 AVSS.n594 17.6946
R2095 AVSS.n551 AVSS.n550 17.6946
R2096 AVSS.n1453 AVSS.n1451 17.6946
R2097 AVSS.n1515 AVSS.n1514 17.6946
R2098 AVSS.n1023 AVSS.n198 17.6946
R2099 AVSS.n844 AVSS.n843 17.6946
R2100 AVSS.n1643 AVSS.t65 17.4005
R2101 AVSS.n1643 AVSS.t56 17.4005
R2102 AVSS.n1610 AVSS.t107 17.4005
R2103 AVSS.n1610 AVSS.t45 17.4005
R2104 AVSS.t83 AVSS.n1177 17.4005
R2105 AVSS.n1177 AVSS.t126 17.4005
R2106 AVSS.t162 AVSS.n1013 17.4005
R2107 AVSS.n1013 AVSS.t41 17.4005
R2108 AVSS.n926 AVSS.t63 17.4005
R2109 AVSS.n926 AVSS.t53 17.4005
R2110 AVSS.n719 AVSS.t31 17.4005
R2111 AVSS.n719 AVSS.t27 17.4005
R2112 AVSS.n656 AVSS.t120 17.4005
R2113 AVSS.n656 AVSS.t115 17.4005
R2114 AVSS.n1060 AVSS.t67 17.4005
R2115 AVSS.n1060 AVSS.t135 17.4005
R2116 AVSS.n1059 AVSS.t72 17.4005
R2117 AVSS.t67 AVSS.n1059 17.4005
R2118 AVSS.t164 AVSS.n240 17.4005
R2119 AVSS.n240 AVSS.t72 17.4005
R2120 AVSS.t89 AVSS.n820 17.4005
R2121 AVSS.n820 AVSS.t12 17.4005
R2122 AVSS.n821 AVSS.t91 17.4005
R2123 AVSS.n821 AVSS.t89 17.4005
R2124 AVSS.n819 AVSS.t38 17.4005
R2125 AVSS.t91 AVSS.n819 17.4005
R2126 AVSS.t118 AVSS.n397 17.4005
R2127 AVSS.n397 AVSS.t112 17.4005
R2128 AVSS.t24 AVSS.n613 17.4005
R2129 AVSS.n613 AVSS.t19 17.4005
R2130 AVSS.t16 AVSS.n449 17.4005
R2131 AVSS.n449 AVSS.t178 17.4005
R2132 AVSS.t80 AVSS.n476 17.4005
R2133 AVSS.n476 AVSS.t74 17.4005
R2134 AVSS.t22 AVSS.n523 17.4005
R2135 AVSS.n523 AVSS.t138 17.4005
R2136 AVSS.n1264 AVSS.t70 17.4005
R2137 AVSS.n1264 AVSS.t151 17.4005
R2138 AVSS.n1198 AVSS.t110 17.4005
R2139 AVSS.n1198 AVSS.t172 17.4005
R2140 AVSS.n1033 AVSS.t155 17.4005
R2141 AVSS.n1033 AVSS.t147 17.4005
R2142 AVSS.n953 AVSS.t167 17.4005
R2143 AVSS.n953 AVSS.t158 17.4005
R2144 AVSS.t133 AVSS.n308 17.4005
R2145 AVSS.n308 AVSS.t9 17.4005
R2146 AVSS.t60 AVSS.n1397 17.4005
R2147 AVSS.n1397 AVSS.t49 17.4005
R2148 AVSS.t104 AVSS.n1384 17.4005
R2149 AVSS.n1384 AVSS.t98 17.4005
R2150 AVSS.t96 AVSS.n1359 17.4005
R2151 AVSS.n1359 AVSS.t93 17.4005
R2152 AVSS.t144 AVSS.n1488 17.4005
R2153 AVSS.n1488 AVSS.t141 17.4005
R2154 AVSS.t169 AVSS.n1328 17.4005
R2155 AVSS.n1328 AVSS.t122 17.4005
R2156 AVSS.n424 AVSS.n422 16.9417
R2157 AVSS.n469 AVSS.n467 16.9417
R2158 AVSS.n1431 AVSS.n1379 16.9417
R2159 AVSS.n1493 AVSS.n1349 16.9417
R2160 AVSS.n1553 AVSS.n1320 16.9417
R2161 AVSS.n875 AVSS.n785 16.9417
R2162 AVSS.n1071 AVSS.n1070 16.9417
R2163 AVSS.n11 AVSS.n1 16.9417
R2164 AVSS.n824 AVSS.n816 16.9417
R2165 AVSS.n372 AVSS.n367 16.5652
R2166 AVSS.n317 AVSS.n310 16.5652
R2167 AVSS.n749 AVSS.n747 16.5652
R2168 AVSS.n996 AVSS.n222 16.5652
R2169 AVSS.n1165 AVSS.n110 16.5652
R2170 AVSS.n78 AVSS.n72 16.5652
R2171 AVSS.n1719 AVSS.n1258 16.5652
R2172 AVSS.n1280 AVSS.n1279 16.5652
R2173 AVSS.n663 AVSS.n662 16.5652
R2174 AVSS.n728 AVSS.n727 16.5652
R2175 AVSS.n741 AVSS.n329 16.5652
R2176 AVSS.n1008 AVSS.n215 16.5652
R2177 AVSS.n1153 AVSS.n1152 16.5652
R2178 AVSS.n1183 AVSS.n66 16.5652
R2179 AVSS.n1596 AVSS.n1575 16.5652
R2180 AVSS.n1627 AVSS.n1626 16.5652
R2181 AVSS.t33 AVSS.n279 16.2348
R2182 AVSS.t59 AVSS.n1290 16.2348
R2183 AVSS.n435 AVSS.n433 16.1887
R2184 AVSS.n486 AVSS.n484 16.1887
R2185 AVSS.n1374 AVSS.n1373 16.1887
R2186 AVSS.n1344 AVSS.n1343 16.1887
R2187 AVSS.n1316 AVSS.n1313 16.1887
R2188 AVSS.n1022 AVSS.n199 16.1887
R2189 AVSS.n842 AVSS.n808 16.1887
R2190 AVSS.n1138 AVSS.t5 15.7275
R2191 AVSS.n605 AVSS.n426 15.4358
R2192 AVSS.n562 AVSS.n471 15.4358
R2193 AVSS.n1438 AVSS.n1378 15.4358
R2194 AVSS.n1500 AVSS.n1348 15.4358
R2195 AVSS.n1667 AVSS.n1666 15.4358
R2196 AVSS.n872 AVSS.n789 15.4358
R2197 AVSS.n176 AVSS.n153 15.4358
R2198 AVSS.n1756 AVSS.n1755 15.4358
R2199 AVSS.n833 AVSS.n831 15.4358
R2200 AVSS.n1162 AVSS.t5 15.2201
R2201 AVSS.n648 AVSS.n362 15.0593
R2202 AVSS.n684 AVSS.n368 15.0593
R2203 AVSS.n763 AVSS.n318 15.0593
R2204 AVSS.n757 AVSS.n325 15.0593
R2205 AVSS.n1170 AVSS.n1168 15.0593
R2206 AVSS.n1194 AVSS.n82 15.0593
R2207 AVSS.n1718 AVSS.n1259 15.0593
R2208 AVSS.n1711 AVSS.n1270 15.0593
R2209 AVSS.n653 AVSS.n652 15.0593
R2210 AVSS.n664 AVSS.n660 15.0593
R2211 AVSS.n729 AVSS.n331 15.0593
R2212 AVSS.n738 AVSS.n737 15.0593
R2213 AVSS.n1174 AVSS.n103 15.0593
R2214 AVSS.n1184 AVSS.n1182 15.0593
R2215 AVSS.n1617 AVSS.n1616 15.0593
R2216 AVSS.n1625 AVSS.n1572 15.0593
R2217 AVSS.n932 AVSS.t33 14.7128
R2218 AVSS.n600 AVSS.n431 14.6829
R2219 AVSS.n556 AVSS.n482 14.6829
R2220 AVSS.n1445 AVSS.n1444 14.6829
R2221 AVSS.n1508 AVSS.n1507 14.6829
R2222 AVSS.n1673 AVSS.n1317 14.6829
R2223 AVSS.n203 AVSS.n202 14.6829
R2224 AVSS.n815 AVSS.n811 14.6829
R2225 AVSS.n604 AVSS.n427 13.9299
R2226 AVSS.n561 AVSS.n472 13.9299
R2227 AVSS.n1440 AVSS.n1439 13.9299
R2228 AVSS.n1502 AVSS.n1501 13.9299
R2229 AVSS.n1318 AVSS.n1315 13.9299
R2230 AVSS.n1046 AVSS.n1045 13.9299
R2231 AVSS.n835 AVSS.n834 13.9299
R2232 AVSS.n370 AVSS.n361 13.5534
R2233 AVSS.n685 AVSS.n370 13.5534
R2234 AVSS.n762 AVSS.n319 13.5534
R2235 AVSS.n758 AVSS.n319 13.5534
R2236 AVSS.n1169 AVSS.n77 13.5534
R2237 AVSS.n1195 AVSS.n77 13.5534
R2238 AVSS.n1269 AVSS.n1268 13.5534
R2239 AVSS.n1712 AVSS.n1269 13.5534
R2240 AVSS.n389 AVSS.n382 13.5534
R2241 AVSS.n659 AVSS.n382 13.5534
R2242 AVSS.n735 AVSS.n733 13.5534
R2243 AVSS.n736 AVSS.n735 13.5534
R2244 AVSS.n1175 AVSS.n101 13.5534
R2245 AVSS.n1181 AVSS.n101 13.5534
R2246 AVSS.n1620 AVSS.n1574 13.5534
R2247 AVSS.n1621 AVSS.n1620 13.5534
R2248 AVSS.n601 AVSS.n427 13.177
R2249 AVSS.n557 AVSS.n472 13.177
R2250 AVSS.n1439 AVSS.n1376 13.177
R2251 AVSS.n1501 AVSS.n1346 13.177
R2252 AVSS.n1674 AVSS.n1318 13.177
R2253 AVSS.n1046 AVSS.n175 13.177
R2254 AVSS.n836 AVSS.n835 13.177
R2255 AVSS.t8 AVSS.n766 12.6835
R2256 AVSS.n601 AVSS.n600 12.424
R2257 AVSS.n557 AVSS.n556 12.424
R2258 AVSS.n1445 AVSS.n1376 12.424
R2259 AVSS.n1508 AVSS.n1346 12.424
R2260 AVSS.n1674 AVSS.n1673 12.424
R2261 AVSS.n202 AVSS.n175 12.424
R2262 AVSS.n836 AVSS.n815 12.424
R2263 AVSS.n648 AVSS.n361 12.0476
R2264 AVSS.n685 AVSS.n684 12.0476
R2265 AVSS.n763 AVSS.n762 12.0476
R2266 AVSS.n758 AVSS.n757 12.0476
R2267 AVSS.n1170 AVSS.n1169 12.0476
R2268 AVSS.n1195 AVSS.n1194 12.0476
R2269 AVSS.n1268 AVSS.n1259 12.0476
R2270 AVSS.n1712 AVSS.n1711 12.0476
R2271 AVSS.n652 AVSS.n389 12.0476
R2272 AVSS.n660 AVSS.n659 12.0476
R2273 AVSS.n733 AVSS.n331 12.0476
R2274 AVSS.n737 AVSS.n736 12.0476
R2275 AVSS.n1175 AVSS.n1174 12.0476
R2276 AVSS.n1182 AVSS.n1181 12.0476
R2277 AVSS.n1617 AVSS.n1574 12.0476
R2278 AVSS.n1621 AVSS.n1572 12.0476
R2279 AVSS.n605 AVSS.n604 11.6711
R2280 AVSS.n562 AVSS.n561 11.6711
R2281 AVSS.n1440 AVSS.n1438 11.6711
R2282 AVSS.n1502 AVSS.n1500 11.6711
R2283 AVSS.n1667 AVSS.n1315 11.6711
R2284 AVSS.n1045 AVSS.n176 11.6711
R2285 AVSS.n834 AVSS.n833 11.6711
R2286 AVSS.n433 AVSS.n431 10.9181
R2287 AVSS.n484 AVSS.n482 10.9181
R2288 AVSS.n1444 AVSS.n1374 10.9181
R2289 AVSS.n1507 AVSS.n1344 10.9181
R2290 AVSS.n1317 AVSS.n1316 10.9181
R2291 AVSS.n203 AVSS.n199 10.9181
R2292 AVSS.n811 AVSS.n808 10.9181
R2293 AVSS.n646 AVSS.n362 10.5417
R2294 AVSS.n372 AVSS.n368 10.5417
R2295 AVSS.n318 AVSS.n317 10.5417
R2296 AVSS.n747 AVSS.n325 10.5417
R2297 AVSS.n1168 AVSS.n110 10.5417
R2298 AVSS.n82 AVSS.n78 10.5417
R2299 AVSS.n1719 AVSS.n1718 10.5417
R2300 AVSS.n1279 AVSS.n1270 10.5417
R2301 AVSS.n653 AVSS.n387 10.5417
R2302 AVSS.n664 AVSS.n663 10.5417
R2303 AVSS.n729 AVSS.n728 10.5417
R2304 AVSS.n738 AVSS.n329 10.5417
R2305 AVSS.n1152 AVSS.n103 10.5417
R2306 AVSS.n1184 AVSS.n1183 10.5417
R2307 AVSS.n1616 AVSS.n1575 10.5417
R2308 AVSS.n1626 AVSS.n1625 10.5417
R2309 AVSS.n426 AVSS.n424 10.1652
R2310 AVSS.n471 AVSS.n469 10.1652
R2311 AVSS.n1379 AVSS.n1378 10.1652
R2312 AVSS.n1349 AVSS.n1348 10.1652
R2313 AVSS.n1666 AVSS.n1320 10.1652
R2314 AVSS.n875 AVSS.n789 10.1652
R2315 AVSS.n1071 AVSS.n153 10.1652
R2316 AVSS.n1756 AVSS.n11 10.1652
R2317 AVSS.n831 AVSS.n816 10.1652
R2318 AVSS.n946 AVSS.t1 9.63961
R2319 AVSS.n595 AVSS.n435 9.41227
R2320 AVSS.n551 AVSS.n486 9.41227
R2321 AVSS.n1451 AVSS.n1373 9.41227
R2322 AVSS.n1514 AVSS.n1343 9.41227
R2323 AVSS.n1023 AVSS.n1022 9.41227
R2324 AVSS.n843 AVSS.n842 9.41227
R2325 AVSS.n686 AVSS.n685 9.3005
R2326 AVSS.n686 AVSS.n368 9.3005
R2327 AVSS.n686 AVSS.n367 9.3005
R2328 AVSS.n686 AVSS.n366 9.3005
R2329 AVSS.n686 AVSS.n365 9.3005
R2330 AVSS.n686 AVSS.n359 9.3005
R2331 AVSS.n687 AVSS.n686 9.3005
R2332 AVSS.n686 AVSS.n363 9.3005
R2333 AVSS.n759 AVSS.n758 9.3005
R2334 AVSS.n325 AVSS.n324 9.3005
R2335 AVSS.n749 AVSS.n748 9.3005
R2336 AVSS.n750 AVSS.n266 9.3005
R2337 AVSS.n951 AVSS.n950 9.3005
R2338 AVSS.n269 AVSS.n267 9.3005
R2339 AVSS.n940 AVSS.n939 9.3005
R2340 AVSS.n942 AVSS.n265 9.3005
R2341 AVSS.n1000 AVSS.n222 9.3005
R2342 AVSS.n1002 AVSS.n1001 9.3005
R2343 AVSS.n190 AVSS.n186 9.3005
R2344 AVSS.n1031 AVSS.n1030 9.3005
R2345 AVSS.n187 AVSS.n183 9.3005
R2346 AVSS.n1036 AVSS.n1035 9.3005
R2347 AVSS.n1196 AVSS.n1195 9.3005
R2348 AVSS.n82 AVSS.n81 9.3005
R2349 AVSS.n74 AVSS.n72 9.3005
R2350 AVSS.n1206 AVSS.n1205 9.3005
R2351 AVSS.n1201 AVSS.n1200 9.3005
R2352 AVSS.n56 AVSS.n55 9.3005
R2353 AVSS.n1234 AVSS.n1233 9.3005
R2354 AVSS.n1236 AVSS.n54 9.3005
R2355 AVSS.n1713 AVSS.n1712 9.3005
R2356 AVSS.n1270 AVSS.n1267 9.3005
R2357 AVSS.n1283 AVSS.n1280 9.3005
R2358 AVSS.n1704 AVSS.n1703 9.3005
R2359 AVSS.n1702 AVSS.n1701 9.3005
R2360 AVSS.n1285 AVSS.n1284 9.3005
R2361 AVSS.n1692 AVSS.n1293 9.3005
R2362 AVSS.n1693 AVSS.n1692 9.3005
R2363 AVSS.n686 AVSS.n362 9.3005
R2364 AVSS.n686 AVSS.n361 9.3005
R2365 AVSS.n703 AVSS.n702 9.3005
R2366 AVSS.n705 AVSS.n342 9.3005
R2367 AVSS.n710 AVSS.n709 9.3005
R2368 AVSS.n706 AVSS.n305 9.3005
R2369 AVSS.n774 AVSS.n773 9.3005
R2370 AVSS.n771 AVSS.n770 9.3005
R2371 AVSS.n320 AVSS.n310 9.3005
R2372 AVSS.n323 AVSS.n318 9.3005
R2373 AVSS.n762 AVSS.n761 9.3005
R2374 AVSS.n955 AVSS.n263 9.3005
R2375 AVSS.n964 AVSS.n963 9.3005
R2376 AVSS.n960 AVSS.n959 9.3005
R2377 AVSS.n229 AVSS.n228 9.3005
R2378 AVSS.n998 AVSS.n997 9.3005
R2379 AVSS.n146 AVSS.n145 9.3005
R2380 AVSS.n1079 AVSS.n1078 9.3005
R2381 AVSS.n144 AVSS.n142 9.3005
R2382 AVSS.n1088 AVSS.n1087 9.3005
R2383 AVSS.n1085 AVSS.n1084 9.3005
R2384 AVSS.n112 AVSS.n111 9.3005
R2385 AVSS.n1166 AVSS.n1165 9.3005
R2386 AVSS.n1168 AVSS.n1167 9.3005
R2387 AVSS.n1169 AVSS.n75 9.3005
R2388 AVSS.n1737 AVSS.n1237 9.3005
R2389 AVSS.n1581 AVSS.n1238 9.3005
R2390 AVSS.n1580 AVSS.n1246 9.3005
R2391 AVSS.n1729 AVSS.n1728 9.3005
R2392 AVSS.n1727 AVSS.n1726 9.3005
R2393 AVSS.n1260 AVSS.n1250 9.3005
R2394 AVSS.n1263 AVSS.n1258 9.3005
R2395 AVSS.n1718 AVSS.n1717 9.3005
R2396 AVSS.n1268 AVSS.n1266 9.3005
R2397 AVSS.n1692 AVSS.n1297 9.3005
R2398 AVSS.n1692 AVSS.n1299 9.3005
R2399 AVSS.n1692 AVSS.n1296 9.3005
R2400 AVSS.n1692 AVSS.n1300 9.3005
R2401 AVSS.n1692 AVSS.n1295 9.3005
R2402 AVSS.n1692 AVSS.n1691 9.3005
R2403 AVSS.n537 AVSS.n536 9.3005
R2404 AVSS.n540 AVSS.n539 9.3005
R2405 AVSS.n496 AVSS.n494 9.3005
R2406 AVSS.n490 AVSS.n489 9.3005
R2407 AVSS.n548 AVSS.n547 9.3005
R2408 AVSS.n550 AVSS.n549 9.3005
R2409 AVSS.n488 AVSS.n486 9.3005
R2410 AVSS.n482 AVSS.n481 9.3005
R2411 AVSS.n558 AVSS.n557 9.3005
R2412 AVSS.n456 AVSS.n451 9.3005
R2413 AVSS.n584 AVSS.n583 9.3005
R2414 AVSS.n446 AVSS.n443 9.3005
R2415 AVSS.n439 AVSS.n438 9.3005
R2416 AVSS.n592 AVSS.n591 9.3005
R2417 AVSS.n594 AVSS.n593 9.3005
R2418 AVSS.n437 AVSS.n435 9.3005
R2419 AVSS.n431 AVSS.n430 9.3005
R2420 AVSS.n602 AVSS.n601 9.3005
R2421 AVSS.n412 AVSS.n410 9.3005
R2422 AVSS.n402 AVSS.n399 9.3005
R2423 AVSS.n637 AVSS.n636 9.3005
R2424 AVSS.n400 AVSS.n396 9.3005
R2425 AVSS.n642 AVSS.n641 9.3005
R2426 AVSS.n645 AVSS.n644 9.3005
R2427 AVSS.n512 AVSS.n510 9.3005
R2428 AVSS.n514 AVSS.n513 9.3005
R2429 AVSS.n511 AVSS.n509 9.3005
R2430 AVSS.n506 AVSS.n505 9.3005
R2431 AVSS.n522 AVSS.n521 9.3005
R2432 AVSS.n529 AVSS.n528 9.3005
R2433 AVSS.n501 AVSS.n497 9.3005
R2434 AVSS.n561 AVSS.n560 9.3005
R2435 AVSS.n480 AVSS.n471 9.3005
R2436 AVSS.n473 AVSS.n467 9.3005
R2437 AVSS.n569 AVSS.n568 9.3005
R2438 AVSS.n571 AVSS.n570 9.3005
R2439 AVSS.n465 AVSS.n463 9.3005
R2440 AVSS.n454 AVSS.n452 9.3005
R2441 AVSS.n579 AVSS.n578 9.3005
R2442 AVSS.n604 AVSS.n603 9.3005
R2443 AVSS.n429 AVSS.n426 9.3005
R2444 AVSS.n422 AVSS.n421 9.3005
R2445 AVSS.n612 AVSS.n611 9.3005
R2446 AVSS.n619 AVSS.n618 9.3005
R2447 AVSS.n414 AVSS.n413 9.3005
R2448 AVSS.n626 AVSS.n625 9.3005
R2449 AVSS.n628 AVSS.n627 9.3005
R2450 AVSS.n1530 AVSS.n1330 9.3005
R2451 AVSS.n1528 AVSS.n1527 9.3005
R2452 AVSS.n1525 AVSS.n1524 9.3005
R2453 AVSS.n1337 AVSS.n1336 9.3005
R2454 AVSS.n1518 AVSS.n1517 9.3005
R2455 AVSS.n1516 AVSS.n1515 9.3005
R2456 AVSS.n1343 AVSS.n1342 9.3005
R2457 AVSS.n1507 AVSS.n1506 9.3005
R2458 AVSS.n1505 AVSS.n1346 9.3005
R2459 AVSS.n1363 AVSS.n1357 9.3005
R2460 AVSS.n1468 AVSS.n1467 9.3005
R2461 AVSS.n1368 AVSS.n1361 9.3005
R2462 AVSS.n1458 AVSS.n1457 9.3005
R2463 AVSS.n1455 AVSS.n1371 9.3005
R2464 AVSS.n1454 AVSS.n1453 9.3005
R2465 AVSS.n1373 AVSS.n1372 9.3005
R2466 AVSS.n1444 AVSS.n1443 9.3005
R2467 AVSS.n1442 AVSS.n1376 9.3005
R2468 AVSS.n1412 AVSS.n1411 9.3005
R2469 AVSS.n1403 AVSS.n1392 9.3005
R2470 AVSS.n1402 AVSS.n1401 9.3005
R2471 AVSS.n1395 AVSS.n1304 9.3005
R2472 AVSS.n1687 AVSS.n1686 9.3005
R2473 AVSS.n1414 AVSS.n1413 9.3005
R2474 AVSS.n1415 AVSS.n1386 9.3005
R2475 AVSS.n1424 AVSS.n1423 9.3005
R2476 AVSS.n1389 AVSS.n1382 9.3005
R2477 AVSS.n1428 AVSS.n1381 9.3005
R2478 AVSS.n1431 AVSS.n1430 9.3005
R2479 AVSS.n1378 AVSS.n1377 9.3005
R2480 AVSS.n1441 AVSS.n1440 9.3005
R2481 AVSS.n1472 AVSS.n1356 9.3005
R2482 AVSS.n1474 AVSS.n1473 9.3005
R2483 AVSS.n1353 AVSS.n1352 9.3005
R2484 AVSS.n1484 AVSS.n1483 9.3005
R2485 AVSS.n1485 AVSS.n1351 9.3005
R2486 AVSS.n1493 AVSS.n1492 9.3005
R2487 AVSS.n1348 AVSS.n1347 9.3005
R2488 AVSS.n1503 AVSS.n1502 9.3005
R2489 AVSS.n1539 AVSS.n1538 9.3005
R2490 AVSS.n1333 AVSS.n1326 9.3005
R2491 AVSS.n1543 AVSS.n1325 9.3005
R2492 AVSS.n1545 AVSS.n1544 9.3005
R2493 AVSS.n1322 AVSS.n1321 9.3005
R2494 AVSS.n1554 AVSS.n1553 9.3005
R2495 AVSS.n1666 AVSS.n1665 9.3005
R2496 AVSS.n1690 AVSS.n1689 9.3005
R2497 AVSS.n834 AVSS.n810 9.3005
R2498 AVSS.n831 AVSS.n830 9.3005
R2499 AVSS.n825 AVSS.n824 9.3005
R2500 AVSS.n826 AVSS.n136 9.3005
R2501 AVSS.n1097 AVSS.n1096 9.3005
R2502 AVSS.n1098 AVSS.n133 9.3005
R2503 AVSS.n1135 AVSS.n1134 9.3005
R2504 AVSS.n1131 AVSS.n1130 9.3005
R2505 AVSS.n1104 AVSS.n1102 9.3005
R2506 AVSS.n837 AVSS.n836 9.3005
R2507 AVSS.n811 AVSS.n809 9.3005
R2508 AVSS.n842 AVSS.n841 9.3005
R2509 AVSS.n845 AVSS.n844 9.3005
R2510 AVSS.n849 AVSS.n848 9.3005
R2511 AVSS.n817 AVSS.n803 9.3005
R2512 AVSS.n854 AVSS.n802 9.3005
R2513 AVSS.n857 AVSS.n856 9.3005
R2514 AVSS.n859 AVSS.n858 9.3005
R2515 AVSS.n870 AVSS.n869 9.3005
R2516 AVSS.n798 AVSS.n796 9.3005
R2517 AVSS.n865 AVSS.n864 9.3005
R2518 AVSS.n899 AVSS.n786 9.3005
R2519 AVSS.n899 AVSS.n788 9.3005
R2520 AVSS.n900 AVSS.n899 9.3005
R2521 AVSS.n899 AVSS.n789 9.3005
R2522 AVSS.n899 AVSS.n785 9.3005
R2523 AVSS.n899 AVSS.n790 9.3005
R2524 AVSS.n899 AVSS.n784 9.3005
R2525 AVSS.n899 AVSS.n791 9.3005
R2526 AVSS.n899 AVSS.n783 9.3005
R2527 AVSS.n899 AVSS.n898 9.3005
R2528 AVSS.n902 AVSS.n287 9.3005
R2529 AVSS.n1748 AVSS.n1747 9.3005
R2530 AVSS.n291 AVSS.n287 9.3005
R2531 AVSS.n1749 AVSS.n1748 9.3005
R2532 AVSS.n908 AVSS.n287 9.3005
R2533 AVSS.n916 AVSS.n910 9.3005
R2534 AVSS.n911 AVSS.n282 9.3005
R2535 AVSS.n929 AVSS.n928 9.3005
R2536 AVSS.n972 AVSS.n257 9.3005
R2537 AVSS.n1045 AVSS.n1044 9.3005
R2538 AVSS.n169 AVSS.n153 9.3005
R2539 AVSS.n1070 AVSS.n1069 9.3005
R2540 AVSS.n167 AVSS.n166 9.3005
R2541 AVSS.n1061 AVSS.n128 9.3005
R2542 AVSS.n1145 AVSS.n1144 9.3005
R2543 AVSS.n1148 AVSS.n119 9.3005
R2544 AVSS.n1158 AVSS.n1157 9.3005
R2545 AVSS.n659 AVSS.n658 9.3005
R2546 AVSS.n665 AVSS.n664 9.3005
R2547 AVSS.n662 AVSS.n380 9.3005
R2548 AVSS.n669 AVSS.n378 9.3005
R2549 AVSS.n672 AVSS.n671 9.3005
R2550 AVSS.n352 AVSS.n351 9.3005
R2551 AVSS.n694 AVSS.n693 9.3005
R2552 AVSS.n696 AVSS.n695 9.3005
R2553 AVSS.n736 AVSS.n330 9.3005
R2554 AVSS.n739 AVSS.n738 9.3005
R2555 AVSS.n741 AVSS.n740 9.3005
R2556 AVSS.n742 AVSS.n286 9.3005
R2557 AVSS.n924 AVSS.n923 9.3005
R2558 AVSS.n921 AVSS.n920 9.3005
R2559 AVSS.n916 AVSS.n915 9.3005
R2560 AVSS.n913 AVSS.n911 9.3005
R2561 AVSS.n1009 AVSS.n1008 9.3005
R2562 AVSS.n1011 AVSS.n213 9.3005
R2563 AVSS.n1016 AVSS.n1015 9.3005
R2564 AVSS.n1020 AVSS.n1019 9.3005
R2565 AVSS.n205 AVSS.n178 9.3005
R2566 AVSS.n1043 AVSS.n1042 9.3005
R2567 AVSS.n1181 AVSS.n1180 9.3005
R2568 AVSS.n1185 AVSS.n1184 9.3005
R2569 AVSS.n96 AVSS.n66 9.3005
R2570 AVSS.n1214 AVSS.n1213 9.3005
R2571 AVSS.n1220 AVSS.n61 9.3005
R2572 AVSS.n1225 AVSS.n1224 9.3005
R2573 AVSS.n1745 AVSS.n1744 9.3005
R2574 AVSS.n1587 AVSS.n47 9.3005
R2575 AVSS.n1622 AVSS.n1621 9.3005
R2576 AVSS.n1625 AVSS.n1624 9.3005
R2577 AVSS.n1627 AVSS.n1571 9.3005
R2578 AVSS.n1630 AVSS.n1629 9.3005
R2579 AVSS.n1632 AVSS.n1631 9.3005
R2580 AVSS.n1634 AVSS.n1566 9.3005
R2581 AVSS.n1641 AVSS.n1640 9.3005
R2582 AVSS.n1638 AVSS.n1568 9.3005
R2583 AVSS.n1675 AVSS.n1317 9.3005
R2584 AVSS.n1675 AVSS.n1674 9.3005
R2585 AVSS.n978 AVSS.n977 9.3005
R2586 AVSS.n239 AVSS.n237 9.3005
R2587 AVSS.n989 AVSS.n988 9.3005
R2588 AVSS.n246 AVSS.n245 9.3005
R2589 AVSS.n242 AVSS.n212 9.3005
R2590 AVSS.n1012 AVSS.n198 9.3005
R2591 AVSS.n1022 AVSS.n1021 9.3005
R2592 AVSS.n204 AVSS.n203 9.3005
R2593 AVSS.n177 AVSS.n175 9.3005
R2594 AVSS.n121 AVSS.n102 9.3005
R2595 AVSS.n1179 AVSS.n91 9.3005
R2596 AVSS.n1188 AVSS.n1187 9.3005
R2597 AVSS.n98 AVSS.n97 9.3005
R2598 AVSS.n1216 AVSS.n1215 9.3005
R2599 AVSS.n1748 AVSS.n43 9.3005
R2600 AVSS.n1219 AVSS.n1218 9.3005
R2601 AVSS.n1675 AVSS.n1315 9.3005
R2602 AVSS.n1675 AVSS.n1313 9.3005
R2603 AVSS.n1677 AVSS.n1676 9.3005
R2604 AVSS.n1661 AVSS.n1312 9.3005
R2605 AVSS.n1660 AVSS.n1659 9.3005
R2606 AVSS.n1556 AVSS.n1555 9.3005
R2607 AVSS.n1646 AVSS.n1645 9.3005
R2608 AVSS.n1565 AVSS.n1563 9.3005
R2609 AVSS.n1612 AVSS.n1574 9.3005
R2610 AVSS.n1616 AVSS.n1615 9.3005
R2611 AVSS.n1596 AVSS.n1576 9.3005
R2612 AVSS.n1602 AVSS.n1601 9.3005
R2613 AVSS.n1604 AVSS.n1578 9.3005
R2614 AVSS.n1608 AVSS.n1607 9.3005
R2615 AVSS.n1594 AVSS.n1577 9.3005
R2616 AVSS.n1592 AVSS.n1591 9.3005
R2617 AVSS.n1589 AVSS.n1588 9.3005
R2618 AVSS.n1176 AVSS.n1175 9.3005
R2619 AVSS.n1156 AVSS.n103 9.3005
R2620 AVSS.n1154 AVSS.n1153 9.3005
R2621 AVSS.n1150 AVSS.n1149 9.3005
R2622 AVSS.n160 AVSS.n127 9.3005
R2623 AVSS.n1065 AVSS.n1064 9.3005
R2624 AVSS.n1068 AVSS.n1067 9.3005
R2625 AVSS.n1054 AVSS.n1053 9.3005
R2626 AVSS.n1057 AVSS.n1056 9.3005
R2627 AVSS.n988 AVSS.n987 9.3005
R2628 AVSS.n985 AVSS.n239 9.3005
R2629 AVSS.n977 AVSS.n248 9.3005
R2630 AVSS.n972 AVSS.n971 9.3005
R2631 AVSS.n928 AVSS.n258 9.3005
R2632 AVSS.n733 AVSS.n732 9.3005
R2633 AVSS.n730 AVSS.n729 9.3005
R2634 AVSS.n727 AVSS.n726 9.3005
R2635 AVSS.n723 AVSS.n722 9.3005
R2636 AVSS.n334 AVSS.n298 9.3005
R2637 AVSS.n781 AVSS.n780 9.3005
R2638 AVSS.n338 AVSS.n336 9.3005
R2639 AVSS.n717 AVSS.n716 9.3005
R2640 AVSS.n698 AVSS.n335 9.3005
R2641 AVSS.n389 AVSS.n388 9.3005
R2642 AVSS.n654 AVSS.n653 9.3005
R2643 AVSS.n1757 AVSS.n5 9.3005
R2644 AVSS.n1757 AVSS.n7 9.3005
R2645 AVSS.n1757 AVSS.n4 9.3005
R2646 AVSS.n1757 AVSS.n8 9.3005
R2647 AVSS.n1757 AVSS.n3 9.3005
R2648 AVSS.n1757 AVSS.n9 9.3005
R2649 AVSS.n1757 AVSS.n2 9.3005
R2650 AVSS.n1757 AVSS.n10 9.3005
R2651 AVSS.n1757 AVSS.n1 9.3005
R2652 AVSS.n1757 AVSS.n1756 9.3005
R2653 AVSS.n1112 AVSS.n12 9.3005
R2654 AVSS.n1116 AVSS.n1115 9.3005
R2655 AVSS.n1109 AVSS.n1107 9.3005
R2656 AVSS.n1122 AVSS.n1121 9.3005
R2657 AVSS.n1124 AVSS.n1123 9.3005
R2658 AVSS.n1191 AVSS.t184 9.13229
R2659 AVSS.n1655 AVSS.t48 9.13229
R2660 AVSS.n678 AVSS.n367 9.03579
R2661 AVSS.n769 AVSS.n310 9.03579
R2662 AVSS.n751 AVSS.n749 9.03579
R2663 AVSS.n1003 AVSS.n222 9.03579
R2664 AVSS.n1165 AVSS.n1164 9.03579
R2665 AVSS.n1207 AVSS.n72 9.03579
R2666 AVSS.n1258 AVSS.n1257 9.03579
R2667 AVSS.n1705 AVSS.n1280 9.03579
R2668 AVSS.n662 AVSS.n661 9.03579
R2669 AVSS.n727 AVSS.n333 9.03579
R2670 AVSS.n743 AVSS.n741 9.03579
R2671 AVSS.n1008 AVSS.n1007 9.03579
R2672 AVSS.n1153 AVSS.n1151 9.03579
R2673 AVSS.n1211 AVSS.n66 9.03579
R2674 AVSS.n1597 AVSS.n1596 9.03579
R2675 AVSS.n1628 AVSS.n1627 9.03579
R2676 AVSS.n610 AVSS.n422 8.65932
R2677 AVSS.n567 AVSS.n467 8.65932
R2678 AVSS.n515 AVSS.n514 8.65932
R2679 AVSS.n1432 AVSS.n1431 8.65932
R2680 AVSS.n1494 AVSS.n1493 8.65932
R2681 AVSS.n1553 AVSS.n1552 8.65932
R2682 AVSS.n877 AVSS.n785 8.65932
R2683 AVSS.n1070 AVSS.n154 8.65932
R2684 AVSS.n34 AVSS.n1 8.65932
R2685 AVSS.n824 AVSS.n823 8.65932
R2686 AVSS.n157 AVSS.t0 8.11764
R2687 AVSS.n645 AVSS.n643 7.90638
R2688 AVSS.n594 AVSS.n436 7.90638
R2689 AVSS.n550 AVSS.n487 7.90638
R2690 AVSS.n1690 AVSS.n1302 7.90638
R2691 AVSS.n1453 AVSS.n1452 7.90638
R2692 AVSS.n1515 AVSS.n1341 7.90638
R2693 AVSS.n241 AVSS.n198 7.90638
R2694 AVSS.n1218 AVSS.n1217 7.90638
R2695 AVSS.n844 AVSS.n805 7.90638
R2696 AVSS.n1108 AVSS.n12 7.90638
R2697 AVSS.n676 AVSS.n366 7.52991
R2698 AVSS.n770 AVSS.n306 7.52991
R2699 AVSS.n750 AVSS.n268 7.52991
R2700 AVSS.n1002 AVSS.n223 7.52991
R2701 AVSS.n1083 AVSS.n112 7.52991
R2702 AVSS.n1206 AVSS.n73 7.52991
R2703 AVSS.n1725 AVSS.n1250 7.52991
R2704 AVSS.n1704 AVSS.n1281 7.52991
R2705 AVSS.n1691 AVSS.n1301 7.52991
R2706 AVSS.n673 AVSS.n378 7.52991
R2707 AVSS.n722 AVSS.n721 7.52991
R2708 AVSS.n742 AVSS.n288 7.52991
R2709 AVSS.n213 AVSS.n211 7.52991
R2710 AVSS.n1150 AVSS.n126 7.52991
R2711 AVSS.n1213 AVSS.n1212 7.52991
R2712 AVSS.n1603 AVSS.n1602 7.52991
R2713 AVSS.n1629 AVSS.n1570 7.52991
R2714 AVSS.n1678 AVSS.n1677 7.52991
R2715 AVSS.n908 AVSS.n907 7.52991
R2716 AVSS.n1750 AVSS.n43 7.52991
R2717 AVSS.n611 AVSS.n418 7.15344
R2718 AVSS.n568 AVSS.n464 7.15344
R2719 AVSS.n509 AVSS.n508 7.15344
R2720 AVSS.n1388 AVSS.n1381 7.15344
R2721 AVSS.n1482 AVSS.n1351 7.15344
R2722 AVSS.n1323 AVSS.n1322 7.15344
R2723 AVSS.n880 AVSS.n790 7.15344
R2724 AVSS.n166 AVSS.n165 7.15344
R2725 AVSS.n32 AVSS.n10 7.15344
R2726 AVSS.n1094 AVSS.n136 7.15344
R2727 AVSS.n642 AVSS.n394 6.4005
R2728 AVSS.n591 AVSS.n590 6.4005
R2729 AVSS.n547 AVSS.n546 6.4005
R2730 AVSS.n1686 AVSS.n1685 6.4005
R2731 AVSS.n1459 AVSS.n1371 6.4005
R2732 AVSS.n1519 AVSS.n1518 6.4005
R2733 AVSS.n244 AVSS.n242 6.4005
R2734 AVSS.n1216 AVSS.n64 6.4005
R2735 AVSS.n850 AVSS.n849 6.4005
R2736 AVSS.n1117 AVSS.n1116 6.4005
R2737 AVSS.n650 AVSS.t15 6.08836
R2738 AVSS.n1753 AVSS.n37 6.08836
R2739 AVSS.n1273 AVSS.t150 6.08836
R2740 AVSS.n365 AVSS.n364 6.02403
R2741 AVSS.n775 AVSS.n774 6.02403
R2742 AVSS.n950 AVSS.n949 6.02403
R2743 AVSS.n997 AVSS.n995 6.02403
R2744 AVSS.n1028 AVSS.n190 6.02403
R2745 AVSS.n1084 AVSS.n143 6.02403
R2746 AVSS.n1200 AVSS.n58 6.02403
R2747 AVSS.n1726 AVSS.n1247 6.02403
R2748 AVSS.n1701 AVSS.n1700 6.02403
R2749 AVSS.n1307 AVSS.n1295 6.02403
R2750 AVSS.n672 AVSS.n379 6.02403
R2751 AVSS.n779 AVSS.n298 6.02403
R2752 AVSS.n923 AVSS.n922 6.02403
R2753 AVSS.n987 AVSS.n986 6.02403
R2754 AVSS.n1017 AVSS.n1016 6.02403
R2755 AVSS.n162 AVSS.n160 6.02403
R2756 AVSS.n1226 AVSS.n61 6.02403
R2757 AVSS.n1606 AVSS.n1604 6.02403
R2758 AVSS.n1633 AVSS.n1632 6.02403
R2759 AVSS.n1658 AVSS.n1312 6.02403
R2760 AVSS.n903 AVSS.n291 6.02403
R2761 AVSS.n1749 AVSS.n44 6.02403
R2762 AVSS.n620 AVSS.n619 5.64756
R2763 AVSS.n572 AVSS.n571 5.64756
R2764 AVSS.n520 AVSS.n506 5.64756
R2765 AVSS.n1422 AVSS.n1389 5.64756
R2766 AVSS.n1483 AVSS.n1481 5.64756
R2767 AVSS.n1546 AVSS.n1545 5.64756
R2768 AVSS.n882 AVSS.n784 5.64756
R2769 AVSS.n910 AVSS.n909 5.64756
R2770 AVSS.n1142 AVSS.n128 5.64756
R2771 AVSS.n29 AVSS.n2 5.64756
R2772 AVSS.n1096 AVSS.n1095 5.64756
R2773 AVSS.t132 AVSS.n301 5.58104
R2774 AVSS.n1228 AVSS.t185 5.58104
R2775 AVSS.n401 AVSS.n400 4.89462
R2776 AVSS.n441 AVSS.n439 4.89462
R2777 AVSS.n492 AVSS.n490 4.89462
R2778 AVSS.n1394 AVSS.n1304 4.89462
R2779 AVSS.n1458 AVSS.n1369 4.89462
R2780 AVSS.n1523 AVSS.n1337 4.89462
R2781 AVSS.n245 AVSS.n238 4.89462
R2782 AVSS.n97 AVSS.n92 4.89462
R2783 AVSS.n853 AVSS.n803 4.89462
R2784 AVSS.n1120 AVSS.n1107 4.89462
R2785 AVSS.n688 AVSS.n359 4.51815
R2786 AVSS.n343 AVSS.n305 4.51815
R2787 AVSS.n935 AVSS.n269 4.51815
R2788 AVSS.n958 AVSS.n229 4.51815
R2789 AVSS.n1030 AVSS.n1029 4.51815
R2790 AVSS.n1089 AVSS.n1088 4.51815
R2791 AVSS.n1231 AVSS.n56 4.51815
R2792 AVSS.n1730 AVSS.n1729 4.51815
R2793 AVSS.n1292 AVSS.n1285 4.51815
R2794 AVSS.n1653 AVSS.n1300 4.51815
R2795 AVSS.n692 AVSS.n352 4.51815
R2796 AVSS.n780 AVSS.n297 4.51815
R2797 AVSS.n921 AVSS.n289 4.51815
R2798 AVSS.n985 AVSS.n984 4.51815
R2799 AVSS.n1019 AVSS.n1018 4.51815
R2800 AVSS.n1066 AVSS.n1065 4.51815
R2801 AVSS.n1225 AVSS.n46 4.51815
R2802 AVSS.n1607 AVSS.n1595 4.51815
R2803 AVSS.n1635 AVSS.n1634 4.51815
R2804 AVSS.n1659 AVSS.n1657 4.51815
R2805 AVSS.n902 AVSS.n901 4.51815
R2806 AVSS.n1747 AVSS.n1746 4.51815
R2807 AVSS.n624 AVSS.n414 4.14168
R2808 AVSS.n463 AVSS.n461 4.14168
R2809 AVSS.n521 AVSS.n502 4.14168
R2810 AVSS.n1423 AVSS.n1387 4.14168
R2811 AVSS.n1354 AVSS.n1353 4.14168
R2812 AVSS.n1332 AVSS.n1325 4.14168
R2813 AVSS.n885 AVSS.n791 4.14168
R2814 AVSS.n930 AVSS.n282 4.14168
R2815 AVSS.n1144 AVSS.n1143 4.14168
R2816 AVSS.n27 AVSS.n9 4.14168
R2817 AVSS.n870 AVSS.n794 4.14168
R2818 AVSS.n1136 AVSS.n133 4.14168
R2819 AVSS.n947 AVSS.n272 3.55175
R2820 AVSS.n945 AVSS.n276 3.55175
R2821 AVSS.n933 AVSS.n932 3.55175
R2822 AVSS.n279 AVSS.n260 3.55175
R2823 AVSS.n981 AVSS.n250 3.55175
R2824 AVSS.n982 AVSS.n231 3.55175
R2825 AVSS.n993 AVSS.n992 3.55175
R2826 AVSS.n234 AVSS.n218 3.55175
R2827 AVSS.n1005 AVSS.n220 3.55175
R2828 AVSS.n219 AVSS.n192 3.55175
R2829 AVSS.n1026 AVSS.n1025 3.55175
R2830 AVSS.n812 AVSS.n195 3.55175
R2831 AVSS.n1039 AVSS.n180 3.55175
R2832 AVSS.n1048 AVSS.n172 3.55175
R2833 AVSS.n1049 AVSS.n148 3.55175
R2834 AVSS.n1074 AVSS.n1073 3.55175
R2835 AVSS.n157 AVSS.n138 3.55175
R2836 AVSS.n1092 AVSS.n1091 3.55175
R2837 AVSS.n1140 AVSS.n130 3.55175
R2838 AVSS.n1139 AVSS.n1138 3.55175
R2839 AVSS.n1162 AVSS.n1161 3.55175
R2840 AVSS.n116 AVSS.n106 3.55175
R2841 AVSS.n1172 AVSS.n108 3.55175
R2842 AVSS.n107 AVSS.n84 3.55175
R2843 AVSS.n1192 AVSS.n1191 3.55175
R2844 AVSS.n87 AVSS.n68 3.55175
R2845 AVSS.n1209 AVSS.n70 3.55175
R2846 AVSS.n69 AVSS.n59 3.55175
R2847 AVSS.n636 AVSS.n635 3.38874
R2848 AVSS.n585 AVSS.n443 3.38874
R2849 AVSS.n541 AVSS.n494 3.38874
R2850 AVSS.n1404 AVSS.n1402 3.38874
R2851 AVSS.n1368 AVSS.n1362 3.38874
R2852 AVSS.n1524 AVSS.n1335 3.38874
R2853 AVSS.n990 AVSS.n989 3.38874
R2854 AVSS.n1189 AVSS.n1188 3.38874
R2855 AVSS.n855 AVSS.n854 3.38874
R2856 AVSS.n1121 AVSS.n1103 3.38874
R2857 AVSS.n70 AVSS.t85 3.04443
R2858 AVSS.n687 AVSS.n360 3.01226
R2859 AVSS.n711 AVSS.n710 3.01226
R2860 AVSS.n943 AVSS.n940 3.01226
R2861 AVSS.n959 AVSS.n264 3.01226
R2862 AVSS.n1037 AVSS.n183 3.01226
R2863 AVSS.n1077 AVSS.n142 3.01226
R2864 AVSS.n1233 AVSS.n1232 3.01226
R2865 AVSS.n1246 AVSS.n1245 3.01226
R2866 AVSS.n1694 AVSS.n1293 3.01226
R2867 AVSS.n1651 AVSS.n1296 3.01226
R2868 AVSS.n693 AVSS.n350 3.01226
R2869 AVSS.n715 AVSS.n338 3.01226
R2870 AVSS.n915 AVSS.n914 3.01226
R2871 AVSS.n970 AVSS.n248 3.01226
R2872 AVSS.n1041 AVSS.n178 3.01226
R2873 AVSS.n1067 AVSS.n159 3.01226
R2874 AVSS.n1744 AVSS.n1743 3.01226
R2875 AVSS.n1594 AVSS.n1593 3.01226
R2876 AVSS.n1640 AVSS.n1639 3.01226
R2877 AVSS.n1564 AVSS.n1556 3.01226
R2878 AVSS.n900 AVSS.n293 3.01226
R2879 AVSS.n38 AVSS.n4 3.01226
R2880 AVSS.n625 AVSS.n411 2.63579
R2881 AVSS.n577 AVSS.n454 2.63579
R2882 AVSS.n530 AVSS.n529 2.63579
R2883 AVSS.n1416 AVSS.n1415 2.63579
R2884 AVSS.n1475 AVSS.n1474 2.63579
R2885 AVSS.n1537 AVSS.n1333 2.63579
R2886 AVSS.n897 AVSS.n783 2.63579
R2887 AVSS.n929 AVSS.n283 2.63579
R2888 AVSS.n1159 AVSS.n119 2.63579
R2889 AVSS.n24 AVSS.n3 2.63579
R2890 AVSS.n799 AVSS.n798 2.63579
R2891 AVSS.n1135 AVSS.n134 2.63579
R2892 AVSS.t30 AVSS.t132 2.53711
R2893 AVSS.t26 AVSS.t8 2.53711
R2894 AVSS.t62 AVSS.t166 2.53711
R2895 AVSS.n967 AVSS.t188 2.53711
R2896 AVSS.t52 AVSS.t157 2.53711
R2897 AVSS.n220 AVSS.t37 2.53711
R2898 AVSS.t161 AVSS.t154 2.53711
R2899 AVSS.t146 AVSS.t40 2.53711
R2900 AVSS.t150 AVSS.t44 2.53711
R2901 AVSS.t82 AVSS.t109 2.02979
R2902 AVSS.t125 AVSS.t171 2.02979
R2903 AVSS.n404 AVSS.n402 1.88285
R2904 AVSS.n584 AVSS.n444 1.88285
R2905 AVSS.n540 AVSS.n495 1.88285
R2906 AVSS.n1403 AVSS.n1393 1.88285
R2907 AVSS.n1467 AVSS.n1466 1.88285
R2908 AVSS.n1529 AVSS.n1528 1.88285
R2909 AVSS.n890 AVSS.n788 1.88285
R2910 AVSS.n254 AVSS.n237 1.88285
R2911 AVSS.n120 AVSS.n91 1.88285
R2912 AVSS.n18 AVSS.n7 1.88285
R2913 AVSS.n856 AVSS.n801 1.88285
R2914 AVSS.n1125 AVSS.n1124 1.88285
R2915 AVSS.t154 AVSS.t3 1.52246
R2916 AVSS.t0 AVSS.t146 1.52246
R2917 AVSS.t184 AVSS.t82 1.52246
R2918 AVSS.t185 AVSS.t125 1.52246
R2919 AVSS.t106 AVSS.t180 1.52246
R2920 AVSS.n1723 AVSS.t106 1.52246
R2921 AVSS.t44 AVSS.t194 1.52246
R2922 AVSS.n363 AVSS.n345 1.50638
R2923 AVSS.n346 AVSS.n342 1.50638
R2924 AVSS.n942 AVSS.n941 1.50638
R2925 AVSS.n965 AVSS.n964 1.50638
R2926 AVSS.n1036 AVSS.n184 1.50638
R2927 AVSS.n1078 AVSS.n1076 1.50638
R2928 AVSS.n1738 AVSS.n54 1.50638
R2929 AVSS.n1736 AVSS.n1238 1.50638
R2930 AVSS.n1693 AVSS.n1294 1.50638
R2931 AVSS.n1560 AVSS.n1299 1.50638
R2932 AVSS.n697 AVSS.n696 1.50638
R2933 AVSS.n716 AVSS.n337 1.50638
R2934 AVSS.n913 AVSS.n912 1.50638
R2935 AVSS.n971 AVSS.n969 1.50638
R2936 AVSS.n1042 AVSS.n170 1.50638
R2937 AVSS.n1055 AVSS.n1054 1.50638
R2938 AVSS.n50 AVSS.n47 1.50638
R2939 AVSS.n1592 AVSS.n1579 1.50638
R2940 AVSS.n1638 AVSS.n1637 1.50638
R2941 AVSS.n1647 AVSS.n1646 1.50638
R2942 AVSS.n629 AVSS.n628 1.12991
R2943 AVSS.n578 AVSS.n453 1.12991
R2944 AVSS.n501 AVSS.n498 1.12991
R2945 AVSS.n1414 AVSS.n1391 1.12991
R2946 AVSS.n1365 AVSS.n1356 1.12991
R2947 AVSS.n1538 AVSS.n1331 1.12991
R2948 AVSS.n898 AVSS.n792 1.12991
R2949 AVSS.n257 AVSS.n253 1.12991
R2950 AVSS.n1158 AVSS.n124 1.12991
R2951 AVSS.n22 AVSS.n8 1.12991
R2952 AVSS.n864 AVSS.n863 1.12991
R2953 AVSS.n1130 AVSS.n1129 1.12991
R2954 AVSS.t18 AVSS.n680 1.01514
R2955 AVSS.t191 AVSS.t30 1.01514
R2956 AVSS.t4 AVSS.t26 1.01514
R2957 AVSS.t1 AVSS.t62 1.01514
R2958 AVSS.t52 AVSS.t188 1.01514
R2959 AVSS.t182 AVSS.t161 1.01514
R2960 AVSS.n1039 AVSS.t3 1.01514
R2961 AVSS.t40 AVSS.t2 1.01514
R2962 AVSS.n1723 AVSS.t69 1.01514
R2963 AVSS.n1586 AVSS.n1585 0.883
R2964 AVSS.n225 AVSS.n224 0.883
R2965 AVSS.n1584 AVSS.n1583 0.88175
R2966 AVSS.n227 AVSS.n226 0.88175
R2967 AVSS.n1583 AVSS.n1582 0.42925
R2968 AVSS.n999 AVSS.n227 0.42925
R2969 AVSS.n1590 AVSS.n1586 0.428
R2970 AVSS.n224 AVSS.n214 0.428
R2971 AVSS.n630 AVSS.n410 0.376971
R2972 AVSS.n457 AVSS.n456 0.376971
R2973 AVSS.n536 AVSS.n535 0.376971
R2974 AVSS.n1411 AVSS.n1410 0.376971
R2975 AVSS.n1366 AVSS.n1363 0.376971
R2976 AVSS.n1531 AVSS.n1530 0.376971
R2977 AVSS.n887 AVSS.n786 0.376971
R2978 AVSS.n979 AVSS.n978 0.376971
R2979 AVSS.n123 AVSS.n121 0.376971
R2980 AVSS.n21 AVSS.n5 0.376971
R2981 AVSS.n860 AVSS.n859 0.376971
R2982 AVSS.n1102 AVSS.n1101 0.376971
R2983 AVSS.n1585 AVSS.n1584 0.3405
R2984 AVSS.n226 AVSS.n225 0.3405
R2985 AVSS.n6 AVSS 0.148784
R2986 AVSS.n899 AVSS.n782 0.105347
R2987 AVSS.n1757 AVSS.n6 0.0999009
R2988 AVSS.n655 AVSS.n384 0.0938044
R2989 AVSS.n381 AVSS 0.0253389
R2990 AVSS.n999 AVSS.n998 0.0247806
R2991 AVSS.n709 AVSS.n705 0.0220827
R2992 AVSS.n761 AVSS.n323 0.0220827
R2993 AVSS.n759 AVSS.n324 0.0220827
R2994 AVSS.n748 AVSS.n324 0.0220827
R2995 AVSS.n748 AVSS.n266 0.0220827
R2996 AVSS.n951 AVSS.n267 0.0220827
R2997 AVSS.n998 AVSS.n228 0.0220827
R2998 AVSS.n1001 AVSS.n1000 0.0220827
R2999 AVSS.n1001 AVSS.n186 0.0220827
R3000 AVSS.n1079 AVSS.n145 0.0220827
R3001 AVSS.n1085 AVSS.n111 0.0220827
R3002 AVSS.n1166 AVSS.n111 0.0220827
R3003 AVSS.n1167 AVSS.n1166 0.0220827
R3004 AVSS.n1167 AVSS.n75 0.0220827
R3005 AVSS.n1234 AVSS.n55 0.0220827
R3006 AVSS.n1237 AVSS.n1236 0.0220827
R3007 AVSS.n1581 AVSS.n1580 0.0220827
R3008 AVSS.n1728 AVSS.n1727 0.0220827
R3009 AVSS.n1713 AVSS.n1267 0.0220827
R3010 AVSS.n1703 AVSS.n1283 0.0220827
R3011 AVSS.n1703 AVSS.n1702 0.0220827
R3012 AVSS.n1702 AVSS.n1284 0.0220827
R3013 AVSS.n939 AVSS.n936 0.0214832
R3014 AVSS.n938 AVSS.n265 0.0214832
R3015 AVSS.n1205 AVSS.n1204 0.0214832
R3016 AVSS.n1202 AVSS.n1201 0.0214832
R3017 AVSS.n1580 AVSS.n1248 0.0211835
R3018 AVSS.n760 AVSS.n759 0.0208837
R3019 AVSS.n858 AVSS.n857 0.0206342
R3020 AVSS.n857 AVSS.n802 0.0206342
R3021 AVSS.n837 AVSS.n810 0.0206342
R3022 AVSS.n1098 AVSS.n1097 0.0206342
R3023 AVSS.n1692 AVSS.n1298 0.0205267
R3024 AVSS.n960 AVSS.n957 0.0199844
R3025 AVSS.n1197 AVSS.n1196 0.0199844
R3026 AVSS.n818 AVSS.n817 0.0197953
R3027 AVSS.n704 AVSS.n703 0.0196847
R3028 AVSS.n703 AVSS.n344 0.0193849
R3029 AVSS.n1080 AVSS.n144 0.0193849
R3030 AVSS.n1087 AVSS.n1082 0.0193849
R3031 AVSS.n1283 AVSS.n1282 0.0193849
R3032 AVSS.n841 AVSS.n840 0.0189564
R3033 AVSS.n838 AVSS.n809 0.0189564
R3034 AVSS.n1134 AVSS.n1099 0.0189564
R3035 AVSS.n1133 AVSS.n1131 0.0189564
R3036 AVSS.n1035 AVSS.n1034 0.0184856
R3037 AVSS.n1717 AVSS.n1716 0.0184856
R3038 AVSS.n1714 AVSS.n1266 0.0184856
R3039 AVSS.n708 AVSS.n706 0.0181859
R3040 AVSS.n773 AVSS.n307 0.0181859
R3041 AVSS.n771 AVSS.n309 0.0169868
R3042 AVSS.n322 AVSS.n320 0.0169868
R3043 AVSS.n1032 AVSS.n1031 0.016687
R3044 AVSS.n1260 AVSS.n1249 0.016687
R3045 AVSS.n1263 AVSS.n1262 0.016687
R3046 AVSS.n686 AVSS.n369 0.0166117
R3047 AVSS.n899 AVSS.n787 0.0165675
R3048 AVSS.n830 AVSS.n822 0.0164396
R3049 AVSS.n826 AVSS.n135 0.0164396
R3050 AVSS.n952 AVSS.n266 0.0163873
R3051 AVSS.n1236 AVSS.n1235 0.0163873
R3052 AVSS.n955 AVSS.n954 0.0151882
R3053 AVSS.n1199 AVSS.n74 0.0151882
R3054 AVSS.n1105 AVSS.n1104 0.0150414
R3055 AVSS.n848 AVSS.n806 0.0139228
R3056 AVSS.n847 AVSS.n845 0.0139228
R3057 AVSS.n956 AVSS.n955 0.0136894
R3058 AVSS.n963 AVSS.n962 0.0136894
R3059 AVSS.n81 AVSS.n76 0.0136894
R3060 AVSS.n80 AVSS.n74 0.0136894
R3061 AVSS.n1086 AVSS.n1085 0.0130899
R3062 AVSS.n845 AVSS.n807 0.0130839
R3063 AVSS.n1104 AVSS.n1100 0.0130839
R3064 AVSS.n869 AVSS.n787 0.0126187
R3065 AVSS AVSS.n0 0.0126187
R3066 AVSS.n1401 AVSS.n1392 0.012516
R3067 AVSS.n1412 AVSS.n1392 0.012516
R3068 AVSS.n1413 AVSS.n1412 0.012516
R3069 AVSS.n1413 AVSS.n1386 0.012516
R3070 AVSS.n1424 AVSS.n1386 0.012516
R3071 AVSS.n1430 AVSS.n1428 0.012516
R3072 AVSS.n1441 AVSS.n1377 0.012516
R3073 AVSS.n1442 AVSS.n1441 0.012516
R3074 AVSS.n1443 AVSS.n1442 0.012516
R3075 AVSS.n1443 AVSS.n1372 0.012516
R3076 AVSS.n1454 AVSS.n1372 0.012516
R3077 AVSS.n1455 AVSS.n1454 0.012516
R3078 AVSS.n1457 AVSS.n1455 0.012516
R3079 AVSS.n1468 AVSS.n1361 0.012516
R3080 AVSS.n1473 AVSS.n1472 0.012516
R3081 AVSS.n1473 AVSS.n1352 0.012516
R3082 AVSS.n1484 AVSS.n1352 0.012516
R3083 AVSS.n1485 AVSS.n1484 0.012516
R3084 AVSS.n1503 AVSS.n1347 0.012516
R3085 AVSS.n1506 AVSS.n1505 0.012516
R3086 AVSS.n1506 AVSS.n1342 0.012516
R3087 AVSS.n1516 AVSS.n1342 0.012516
R3088 AVSS.n1517 AVSS.n1516 0.012516
R3089 AVSS.n1517 AVSS.n1336 0.012516
R3090 AVSS.n1525 AVSS.n1336 0.012516
R3091 AVSS.n1527 AVSS.n1525 0.012516
R3092 AVSS.n1539 AVSS.n1330 0.012516
R3093 AVSS.n1544 AVSS.n1543 0.012516
R3094 AVSS.n1544 AVSS.n1321 0.012516
R3095 AVSS.n1554 AVSS.n1321 0.012516
R3096 AVSS.n1665 AVSS.n1554 0.012516
R3097 AVSS.n1031 AVSS.n189 0.0121906
R3098 AVSS.n187 AVSS.n185 0.0121906
R3099 AVSS.n1265 AVSS.n1263 0.0121906
R3100 AVSS.n1688 AVSS.n1687 0.0120154
R3101 AVSS.n1395 AVSS.n1303 0.0120154
R3102 AVSS.n1401 AVSS.n1400 0.0120154
R3103 AVSS.n772 AVSS.n771 0.0118909
R3104 AVSS.n1665 AVSS.n1664 0.0116816
R3105 AVSS.n1582 AVSS.n1237 0.0112914
R3106 AVSS.n1582 AVSS.n1581 0.0112914
R3107 AVSS.n773 AVSS.n772 0.0106918
R3108 AVSS.n1469 AVSS.n1357 0.0106802
R3109 AVSS.n1472 AVSS.n1471 0.0106802
R3110 AVSS.n830 AVSS.n829 0.0105671
R3111 AVSS.n829 AVSS.n825 0.0105671
R3112 AVSS.n827 AVSS.n825 0.0105671
R3113 AVSS.n827 AVSS.n826 0.0105671
R3114 AVSS.n189 AVSS.n187 0.0103921
R3115 AVSS.n1035 AVSS.n185 0.0103921
R3116 AVSS.n1717 AVSS.n1265 0.0103921
R3117 AVSS.n858 AVSS.n797 0.0103432
R3118 AVSS.n1123 AVSS.n1122 0.0103039
R3119 AVSS.n637 AVSS.n399 0.010167
R3120 AVSS.n412 AVSS.n399 0.010167
R3121 AVSS.n627 AVSS.n412 0.010167
R3122 AVSS.n627 AVSS.n626 0.010167
R3123 AVSS.n626 AVSS.n413 0.010167
R3124 AVSS.n612 AVSS.n421 0.010167
R3125 AVSS.n603 AVSS.n429 0.010167
R3126 AVSS.n603 AVSS.n602 0.010167
R3127 AVSS.n602 AVSS.n430 0.010167
R3128 AVSS.n437 AVSS.n430 0.010167
R3129 AVSS.n593 AVSS.n437 0.010167
R3130 AVSS.n593 AVSS.n592 0.010167
R3131 AVSS.n592 AVSS.n438 0.010167
R3132 AVSS.n583 AVSS.n446 0.010167
R3133 AVSS.n579 AVSS.n452 0.010167
R3134 AVSS.n465 AVSS.n452 0.010167
R3135 AVSS.n570 AVSS.n465 0.010167
R3136 AVSS.n570 AVSS.n569 0.010167
R3137 AVSS.n560 AVSS.n480 0.010167
R3138 AVSS.n558 AVSS.n481 0.010167
R3139 AVSS.n488 AVSS.n481 0.010167
R3140 AVSS.n549 AVSS.n488 0.010167
R3141 AVSS.n549 AVSS.n548 0.010167
R3142 AVSS.n548 AVSS.n489 0.010167
R3143 AVSS.n496 AVSS.n489 0.010167
R3144 AVSS.n539 AVSS.n496 0.010167
R3145 AVSS.n537 AVSS.n497 0.010167
R3146 AVSS.n522 AVSS.n505 0.010167
R3147 AVSS.n511 AVSS.n505 0.010167
R3148 AVSS.n513 AVSS.n511 0.010167
R3149 AVSS.n513 AVSS.n512 0.010167
R3150 AVSS.n641 AVSS.n344 0.00976423
R3151 AVSS.n640 AVSS.n396 0.00976423
R3152 AVSS.n638 AVSS.n637 0.00976423
R3153 AVSS.n868 AVSS.n796 0.00975926
R3154 AVSS.n866 AVSS.n865 0.00975926
R3155 AVSS.n1109 AVSS.n1106 0.00975926
R3156 AVSS.n1429 AVSS.n1377 0.00967891
R3157 AVSS.n512 AVSS.n381 0.0094957
R3158 AVSS.n1087 AVSS.n1086 0.00949281
R3159 AVSS.n1486 AVSS.n1485 0.00901135
R3160 AVSS.n1492 AVSS.n1491 0.00901135
R3161 AVSS.n1540 AVSS.n1326 0.00901135
R3162 AVSS.n1543 AVSS.n1542 0.00901135
R3163 AVSS.n963 AVSS.n956 0.00889329
R3164 AVSS.n962 AVSS.n960 0.00889329
R3165 AVSS.n1196 AVSS.n76 0.00889329
R3166 AVSS.n81 AVSS.n80 0.00889329
R3167 AVSS.n580 AVSS.n579 0.00869012
R3168 AVSS.n1688 AVSS.n1284 0.00859352
R3169 AVSS.n1676 AVSS.n1675 0.00831842
R3170 AVSS.n1505 AVSS.n1504 0.0081769
R3171 AVSS.n1527 AVSS.n1526 0.0081769
R3172 AVSS.n841 AVSS.n807 0.00805034
R3173 AVSS.n1131 AVSS.n1100 0.00805034
R3174 AVSS.n429 AVSS.n428 0.00788453
R3175 AVSS.n1689 AVSS.n1298 0.00784312
R3176 AVSS.n1425 AVSS.n1424 0.00750935
R3177 AVSS.n1427 AVSS.n1382 0.00750935
R3178 AVSS.n954 AVSS.n265 0.00739448
R3179 AVSS.n1205 AVSS.n1199 0.00739448
R3180 AVSS.n569 AVSS.n466 0.00734748
R3181 AVSS.n527 AVSS.n522 0.00734748
R3182 AVSS.n817 AVSS.n806 0.00721141
R3183 AVSS.n848 AVSS.n847 0.00721141
R3184 AVSS.n1115 AVSS.n1110 0.00689978
R3185 AVSS.n1114 AVSS.n1112 0.00689978
R3186 AVSS.n1112 AVSS.n0 0.00676362
R3187 AVSS.n559 AVSS.n558 0.00667615
R3188 AVSS.n539 AVSS.n538 0.00667615
R3189 AVSS.n1457 AVSS.n1456 0.00650801
R3190 AVSS.n1456 AVSS.n1361 0.00650801
R3191 AVSS.n644 AVSS.n369 0.00640763
R3192 AVSS.n952 AVSS.n951 0.00619544
R3193 AVSS.n1235 AVSS.n1234 0.00619544
R3194 AVSS.n419 AVSS.n413 0.0061391
R3195 AVSS.n1032 AVSS.n186 0.00589568
R3196 AVSS.n1727 AVSS.n1249 0.00589568
R3197 AVSS.n1262 AVSS.n1260 0.00589568
R3198 AVSS.n320 AVSS.n309 0.00559592
R3199 AVSS.n323 AVSS.n322 0.00559592
R3200 AVSS.n1425 AVSS.n1382 0.00550668
R3201 AVSS.n1428 AVSS.n1427 0.00550668
R3202 AVSS.n617 AVSS.n616 0.00533351
R3203 AVSS.n445 AVSS.n438 0.00533351
R3204 AVSS.n446 AVSS.n445 0.00533351
R3205 AVSS.n582 AVSS.n448 0.00533351
R3206 AVSS.n479 AVSS.n474 0.00533351
R3207 AVSS.n525 AVSS.n503 0.00533351
R3208 AVSS.n1000 AVSS.n999 0.0049964
R3209 AVSS.n1504 AVSS.n1503 0.00483912
R3210 AVSS.n1526 AVSS.n1330 0.00483912
R3211 AVSS.n822 AVSS.n810 0.00469463
R3212 AVSS.n1097 AVSS.n135 0.00469463
R3213 AVSS.n618 AVSS.n419 0.00452793
R3214 AVSS.n616 AVSS.n612 0.00452793
R3215 AVSS AVSS.n1757 0.0044488
R3216 AVSS.n709 AVSS.n708 0.00439688
R3217 AVSS.n706 AVSS.n307 0.00439688
R3218 AVSS.n655 AVSS.n654 0.0041486
R3219 AVSS.n1034 AVSS.n145 0.00409712
R3220 AVSS.n1716 AVSS.n1266 0.00409712
R3221 AVSS.n1714 AVSS.n1713 0.00409712
R3222 AVSS.n1492 AVSS.n1486 0.00400467
R3223 AVSS.n1491 AVSS.n1347 0.00400467
R3224 AVSS.n1540 AVSS.n1539 0.00400467
R3225 AVSS.n1542 AVSS.n1326 0.00400467
R3226 AVSS.n560 AVSS.n559 0.00399087
R3227 AVSS.n538 AVSS.n537 0.00399087
R3228 AVSS.n671 AVSS.n669 0.00391168
R3229 AVSS.n694 AVSS.n351 0.00391168
R3230 AVSS.n695 AVSS.n694 0.00391168
R3231 AVSS.n695 AVSS.n335 0.00391168
R3232 AVSS.n717 AVSS.n336 0.00391168
R3233 AVSS.n732 AVSS.n330 0.00391168
R3234 AVSS.n739 AVSS.n330 0.00391168
R3235 AVSS.n740 AVSS.n739 0.00391168
R3236 AVSS.n740 AVSS.n286 0.00391168
R3237 AVSS.n916 AVSS.n911 0.00391168
R3238 AVSS.n988 AVSS.n239 0.00391168
R3239 AVSS.n1589 AVSS.n1587 0.00391168
R3240 AVSS.n1591 AVSS.n1577 0.00391168
R3241 AVSS.n1608 AVSS.n1578 0.00391168
R3242 AVSS.n1624 AVSS.n1622 0.00391168
R3243 AVSS.n1630 AVSS.n1571 0.00391168
R3244 AVSS.n1631 AVSS.n1630 0.00391168
R3245 AVSS.n1631 AVSS.n1566 0.00391168
R3246 AVSS.n1641 AVSS.n1568 0.00391168
R3247 AVSS.n1645 AVSS.n1565 0.00391168
R3248 AVSS.n865 AVSS.n797 0.00390414
R3249 AVSS.n1110 AVSS.n1109 0.00390414
R3250 AVSS.n1115 AVSS.n1114 0.00390414
R3251 AVSS.n731 AVSS.n730 0.00386429
R3252 AVSS.n451 AVSS.n448 0.00385661
R3253 AVSS.n247 AVSS.n246 0.00376952
R3254 AVSS.n1623 AVSS.n1571 0.00372214
R3255 AVSS.n334 AVSS.n296 0.0035326
R3256 AVSS.n1609 AVSS.n1577 0.0035326
R3257 AVSS.n1661 AVSS.n1314 0.00348522
R3258 AVSS.n290 AVSS.n287 0.00334306
R3259 AVSS.n977 AVSS.n976 0.00334306
R3260 AVSS.n1430 AVSS.n1429 0.00333712
R3261 AVSS.n473 AVSS.n466 0.00331955
R3262 AVSS.n480 AVSS.n479 0.00331955
R3263 AVSS.n525 AVSS.n497 0.00331955
R3264 AVSS.n528 AVSS.n527 0.00331955
R3265 AVSS.n718 AVSS.n335 0.00329568
R3266 AVSS.n1601 AVSS.n1598 0.00329568
R3267 AVSS.n1600 AVSS.n1576 0.00329568
R3268 AVSS.n666 AVSS.n665 0.00324829
R3269 AVSS.n668 AVSS.n380 0.00324829
R3270 AVSS.n1123 AVSS.n1105 0.00322331
R3271 AVSS.n1587 AVSS.n45 0.00320091
R3272 AVSS.n1080 AVSS.n1079 0.00319784
R3273 AVSS.n1082 AVSS.n144 0.00319784
R3274 AVSS.n1282 AVSS.n1267 0.00319784
R3275 AVSS.n388 AVSS.n386 0.00315353
R3276 AVSS.n658 AVSS.n383 0.00315353
R3277 AVSS.n920 AVSS.n919 0.00310614
R3278 AVSS.n1615 AVSS.n1614 0.00310614
R3279 AVSS.n928 AVSS.n927 0.00305876
R3280 AVSS.n1642 AVSS.n1566 0.0029166
R3281 AVSS.n1644 AVSS.n1555 0.0029166
R3282 AVSS.n705 AVSS.n704 0.00289808
R3283 AVSS.n725 AVSS.n723 0.00286922
R3284 AVSS.n726 AVSS.n332 0.00286922
R3285 AVSS.n1573 AVSS.n6 0.00282183
R3286 AVSS.n428 AVSS.n421 0.00278249
R3287 AVSS.n925 AVSS.n286 0.00277445
R3288 AVSS.n1009 AVSS.n212 0.00277445
R3289 AVSS.n1012 AVSS.n1011 0.00277445
R3290 AVSS.n1044 AVSS.n1043 0.00277445
R3291 AVSS.n1057 AVSS.n169 0.00277445
R3292 AVSS.n1145 AVSS.n127 0.00277445
R3293 AVSS.n1149 AVSS.n1148 0.00277445
R3294 AVSS.n1157 AVSS.n1154 0.00277445
R3295 AVSS.n1219 AVSS.n63 0.00272707
R3296 AVSS.n1567 AVSS.n1565 0.00270571
R3297 AVSS.n1568 AVSS.n1567 0.00270571
R3298 AVSS.n1155 AVSS.n102 0.0026323
R3299 AVSS.n1179 AVSS.n1178 0.0026323
R3300 AVSS.n957 AVSS.n228 0.00259832
R3301 AVSS.n1197 AVSS.n75 0.00259832
R3302 AVSS.n95 AVSS.n65 0.00258491
R3303 AVSS.n1223 AVSS.n62 0.00258491
R3304 AVSS.n723 AVSS.n720 0.00253753
R3305 AVSS.n474 AVSS.n473 0.00251396
R3306 AVSS.n528 AVSS.n503 0.00251396
R3307 AVSS.n1664 AVSS.n1555 0.00249014
R3308 AVSS.n1662 AVSS.n1660 0.00249014
R3309 AVSS.n782 AVSS.n781 0.00244276
R3310 AVSS.n1224 AVSS 0.00234799
R3311 AVSS.n1469 AVSS.n1468 0.00233578
R3312 AVSS.n1471 AVSS.n1357 0.00233578
R3313 AVSS.n1615 AVSS.n1611 0.00230061
R3314 AVSS.n658 AVSS.n657 0.00225322
R3315 AVSS.n1069 AVSS.n155 0.00220584
R3316 AVSS.n167 AVSS.n164 0.00220584
R3317 AVSS.n1590 AVSS.n1589 0.00220584
R3318 AVSS.n1591 AVSS.n1590 0.00220584
R3319 AVSS.n840 AVSS.n809 0.00217785
R3320 AVSS.n838 AVSS.n837 0.00217785
R3321 AVSS.n1099 AVSS.n1098 0.00217785
R3322 AVSS.n1134 AVSS.n1133 0.00217785
R3323 AVSS.n973 AVSS.n256 0.00215845
R3324 AVSS AVSS.n351 0.00211107
R3325 AVSS.n1020 AVSS.n210 0.00211107
R3326 AVSS.n208 AVSS.n205 0.00211107
R3327 AVSS.n1611 AVSS.n1576 0.00211107
R3328 AVSS.n973 AVSS.n972 0.00206368
R3329 AVSS.n977 AVSS.n975 0.00206368
R3330 AVSS.n583 AVSS.n582 0.00197691
R3331 AVSS.n580 AVSS.n451 0.00197691
R3332 AVSS.n670 AVSS 0.00196892
R3333 AVSS.n1664 AVSS.n1660 0.00192153
R3334 AVSS.n1662 AVSS.n1661 0.00192153
R3335 AVSS.n720 AVSS.n334 0.00187415
R3336 AVSS.n1748 AVSS 0.00187415
R3337 AVSS.n1021 AVSS.n200 0.00177938
R3338 AVSS.n761 AVSS.n760 0.00169904
R3339 AVSS.n972 AVSS.n255 0.00168461
R3340 AVSS.n1064 AVSS.n1063 0.00168461
R3341 AVSS.n665 AVSS.n381 0.00163723
R3342 AVSS.n925 AVSS.n924 0.00163723
R3343 AVSS.n1011 AVSS.n212 0.00163723
R3344 AVSS.n1015 AVSS.n1012 0.00163723
R3345 AVSS.n1021 AVSS.n1020 0.00163723
R3346 AVSS.n205 AVSS.n204 0.00163723
R3347 AVSS.n1043 AVSS.n177 0.00163723
R3348 AVSS.n1053 AVSS.n169 0.00163723
R3349 AVSS.n1069 AVSS.n1068 0.00163723
R3350 AVSS.n1064 AVSS.n167 0.00163723
R3351 AVSS.n1061 AVSS.n127 0.00163723
R3352 AVSS.n1157 AVSS.n1156 0.00163723
R3353 AVSS.n1176 AVSS.n102 0.00163723
R3354 AVSS.n1180 AVSS.n1179 0.00163723
R3355 AVSS.n1180 AVSS.n93 0.00163723
R3356 AVSS.n1187 AVSS.n93 0.00163723
R3357 AVSS.n1185 AVSS.n100 0.00163723
R3358 AVSS.n100 AVSS.n98 0.00163723
R3359 AVSS.n98 AVSS.n96 0.00163723
R3360 AVSS.n1215 AVSS.n1214 0.00163723
R3361 AVSS.n782 AVSS.n294 0.00158984
R3362 AVSS.n726 AVSS.n725 0.00154246
R3363 AVSS.n730 AVSS.n332 0.00154246
R3364 AVSS.n1220 AVSS.n62 0.00154246
R3365 AVSS.n1642 AVSS.n1641 0.00149507
R3366 AVSS.n1645 AVSS.n1644 0.00149507
R3367 AVSS.n1186 AVSS.n1185 0.00144769
R3368 AVSS.n1728 AVSS.n1248 0.00139928
R3369 AVSS.n1149 AVSS.n1147 0.00135292
R3370 AVSS.n1154 AVSS.n125 0.00135292
R3371 AVSS.n1221 AVSS.n1219 0.00135292
R3372 AVSS.n818 AVSS.n802 0.00133893
R3373 AVSS.n618 AVSS.n617 0.00130559
R3374 AVSS.n1614 AVSS.n1612 0.00130553
R3375 AVSS.n1622 AVSS.n1573 0.00130553
R3376 AVSS.n654 AVSS.n386 0.00125815
R3377 AVSS.n388 AVSS.n383 0.00125815
R3378 AVSS.n1009 AVSS.n214 0.00121077
R3379 AVSS.n1062 AVSS.n1061 0.00121077
R3380 AVSS.n1745 AVSS.n45 0.00121077
R3381 AVSS.n666 AVSS.n380 0.00116338
R3382 AVSS.n669 AVSS.n668 0.00116338
R3383 AVSS.n919 AVSS.n918 0.00116338
R3384 AVSS.n927 AVSS.n285 0.00116338
R3385 AVSS.n975 AVSS.n255 0.00116338
R3386 AVSS.n718 AVSS.n717 0.001116
R3387 AVSS.n1015 AVSS.n1014 0.001116
R3388 AVSS.n1598 AVSS.n1578 0.001116
R3389 AVSS.n1601 AVSS.n1600 0.001116
R3390 AVSS.n936 AVSS.n267 0.00109952
R3391 AVSS.n939 AVSS.n938 0.00109952
R3392 AVSS.n1204 AVSS.n1201 0.00109952
R3393 AVSS.n1202 AVSS.n55 0.00109952
R3394 AVSS.n976 AVSS.n239 0.00106861
R3395 AVSS.n869 AVSS.n868 0.00104466
R3396 AVSS.n866 AVSS.n796 0.00104466
R3397 AVSS.n1122 AVSS.n1106 0.00104466
R3398 AVSS.n657 AVSS.n381 0.00102123
R3399 AVSS.n1689 AVSS.n1688 0.00100067
R3400 AVSS.n1687 AVSS.n1303 0.00100067
R3401 AVSS.n1400 AVSS.n1395 0.00100067
R3402 AVSS.n924 AVSS.n287 0.000926459
R3403 AVSS.n246 AVSS.n214 0.000926459
R3404 AVSS.n1058 AVSS.n1057 0.000926459
R3405 AVSS.n1676 AVSS.n1314 0.000926459
R3406 AVSS.n644 AVSS.n344 0.000902793
R3407 AVSS.n641 AVSS.n640 0.000902793
R3408 AVSS.n638 AVSS.n396 0.000902793
R3409 AVSS.n336 AVSS.n294 0.000879075
R3410 AVSS.n781 AVSS.n296 0.000879075
R3411 AVSS.n1014 AVSS.n200 0.000879075
R3412 AVSS.n210 AVSS.n201 0.000879075
R3413 AVSS.n208 AVSS.n207 0.000879075
R3414 AVSS.n1058 AVSS.n168 0.000879075
R3415 AVSS.n1052 AVSS.n155 0.000879075
R3416 AVSS.n164 AVSS.n156 0.000879075
R3417 AVSS.n1063 AVSS.n1062 0.000879075
R3418 AVSS.n1609 AVSS.n1608 0.000879075
R3419 AVSS.n671 AVSS.n670 0.000831691
R3420 AVSS.n1044 AVSS.n168 0.000831691
R3421 AVSS.n204 AVSS.n201 0.000784306
R3422 AVSS.n207 AVSS.n177 0.000784306
R3423 AVSS.n1147 AVSS.n1145 0.000784306
R3424 AVSS.n1148 AVSS.n125 0.000784306
R3425 AVSS.n1221 AVSS.n1220 0.000784306
R3426 AVSS.n1224 AVSS.n1223 0.000784306
R3427 AVSS.n1612 AVSS.n6 0.000784306
R3428 AVSS.n911 AVSS.n285 0.000689538
R3429 AVSS.n928 AVSS.n256 0.000689538
R3430 AVSS.n1053 AVSS.n1052 0.000689538
R3431 AVSS.n1068 AVSS.n156 0.000689538
R3432 AVSS.n1187 AVSS.n1186 0.000689538
R3433 AVSS.n1748 AVSS.n1745 0.000689538
R3434 AVSS.n1624 AVSS.n1623 0.000689538
R3435 AVSS.n920 AVSS.n290 0.000642153
R3436 AVSS.n918 AVSS.n916 0.000642153
R3437 AVSS.n988 AVSS.n247 0.000642153
R3438 AVSS.n1156 AVSS.n1155 0.000642153
R3439 AVSS.n1178 AVSS.n1176 0.000642153
R3440 AVSS.n1215 AVSS.n65 0.000642153
R3441 AVSS.n732 AVSS.n731 0.000547384
R3442 AVSS.n96 AVSS.n95 0.000547384
R3443 AVSS.n1214 AVSS.n63 0.000547384
R3444 IREF.n5 IREF.t12 114.496
R3445 IREF.n25 IREF.t10 114.493
R3446 IREF.n52 IREF.t14 114.466
R3447 IREF.n79 IREF.t18 114.466
R3448 IREF.n27 IREF.t20 103.459
R3449 IREF.n20 IREF.t11 103.459
R3450 IREF.n12 IREF.t16 103.459
R3451 IREF.n7 IREF.t13 103.459
R3452 IREF.n36 IREF.t4 103.459
R3453 IREF.n44 IREF.t21 103.459
R3454 IREF.n68 IREF.t8 103.459
R3455 IREF.n60 IREF.t17 103.459
R3456 IREF.n54 IREF.t0 103.459
R3457 IREF.n106 IREF.t24 103.459
R3458 IREF.n113 IREF.t2 103.459
R3459 IREF.n130 IREF.t23 103.459
R3460 IREF.n122 IREF.t6 103.459
R3461 IREF.n94 IREF.t15 103.459
R3462 IREF.n86 IREF.t22 103.459
R3463 IREF.n81 IREF.t19 103.459
R3464 IREF.n70 IREF.t9 87.4858
R3465 IREF.n34 IREF.t5 87.4836
R3466 IREF.n56 IREF.t1 87.4823
R3467 IREF.n118 IREF.t3 87.0905
R3468 IREF.n119 IREF.t7 87.0895
R3469 IREF.n28 IREF.n27 21.9607
R3470 IREF.n27 IREF.n26 21.9607
R3471 IREF.n20 IREF.n19 21.9607
R3472 IREF.n21 IREF.n20 21.9607
R3473 IREF.n12 IREF.n11 21.9607
R3474 IREF.n13 IREF.n12 21.9607
R3475 IREF.n7 IREF.n6 21.9607
R3476 IREF.n8 IREF.n7 21.9607
R3477 IREF.n36 IREF.n35 21.9607
R3478 IREF.n37 IREF.n36 21.9607
R3479 IREF.n45 IREF.n44 21.9607
R3480 IREF.n44 IREF.n43 21.9607
R3481 IREF.n68 IREF.n67 21.9607
R3482 IREF.n69 IREF.n68 21.9607
R3483 IREF.n60 IREF.n59 21.9607
R3484 IREF.n61 IREF.n60 21.9607
R3485 IREF.n54 IREF.n53 21.9607
R3486 IREF.n55 IREF.n54 21.9607
R3487 IREF.n106 IREF.n104 21.9607
R3488 IREF.n107 IREF.n106 21.9607
R3489 IREF.n113 IREF.n102 21.9607
R3490 IREF.n114 IREF.n113 21.9607
R3491 IREF.n130 IREF.n129 21.9607
R3492 IREF.n131 IREF.n130 21.9607
R3493 IREF.n122 IREF.n121 21.9607
R3494 IREF.n123 IREF.n122 21.9607
R3495 IREF.n94 IREF.n93 21.9607
R3496 IREF.n95 IREF.n94 21.9607
R3497 IREF.n86 IREF.n85 21.9607
R3498 IREF.n87 IREF.n86 21.9607
R3499 IREF.n81 IREF.n80 21.9607
R3500 IREF.n82 IREF.n81 21.9607
R3501 IREF.n119 IREF.n118 6.73278
R3502 IREF.n39 IREF.n34 4.61479
R3503 IREF.n117 IREF.n116 4.61479
R3504 IREF.n11 IREF.n10 4.51012
R3505 IREF.n9 IREF.n8 4.51012
R3506 IREF.n22 IREF.n21 4.50915
R3507 IREF.n132 IREF.n131 4.50819
R3508 IREF.n107 IREF.n105 4.50723
R3509 IREF.n85 IREF.n84 4.50539
R3510 IREF.n29 IREF.n28 4.50531
R3511 IREF.n59 IREF.n58 4.50496
R3512 IREF.n96 IREF.n95 4.50406
R3513 IREF.n83 IREF.n82 4.50361
R3514 IREF.n46 IREF.n45 4.50273
R3515 IREF.n24 IREF.n23 4.5005
R3516 IREF.n4 IREF.n3 4.5005
R3517 IREF.n1 IREF.n0 4.5005
R3518 IREF.n18 IREF.n17 4.5005
R3519 IREF.n16 IREF.n2 4.5005
R3520 IREF.n15 IREF.n14 4.5005
R3521 IREF.n39 IREF.n38 4.5005
R3522 IREF.n40 IREF.n33 4.5005
R3523 IREF.n42 IREF.n41 4.5005
R3524 IREF.n32 IREF.n31 4.5005
R3525 IREF.n57 IREF.n56 4.5005
R3526 IREF.n51 IREF.n50 4.5005
R3527 IREF.n71 IREF.n70 4.5005
R3528 IREF.n48 IREF.n47 4.5005
R3529 IREF.n66 IREF.n65 4.5005
R3530 IREF.n64 IREF.n49 4.5005
R3531 IREF.n63 IREF.n62 4.5005
R3532 IREF.n109 IREF.n108 4.5005
R3533 IREF.n111 IREF.n110 4.5005
R3534 IREF.n112 IREF.n103 4.5005
R3535 IREF.n116 IREF.n115 4.5005
R3536 IREF.n99 IREF.n98 4.5005
R3537 IREF.n128 IREF.n127 4.5005
R3538 IREF.n126 IREF.n100 4.5005
R3539 IREF.n125 IREF.n124 4.5005
R3540 IREF.n120 IREF.n101 4.5005
R3541 IREF.n78 IREF.n77 4.5005
R3542 IREF.n75 IREF.n74 4.5005
R3543 IREF.n92 IREF.n91 4.5005
R3544 IREF.n90 IREF.n76 4.5005
R3545 IREF.n89 IREF.n88 4.5005
R3546 IREF.n105 IREF.n101 2.4255
R3547 IREF.n84 IREF.n83 2.4255
R3548 IREF.n10 IREF.n9 2.42193
R3549 IREF.n58 IREF.n57 2.42193
R3550 IREF.n30 IREF.n22 1.89417
R3551 IREF.n72 IREF.n71 1.89381
R3552 IREF.n133 IREF.n132 1.46695
R3553 IREF.n97 IREF.n96 1.4656
R3554 IREF.n79 IREF.n77 1.34987
R3555 IREF.n52 IREF.n50 1.34936
R3556 IREF.n25 IREF.n23 1.33436
R3557 IREF.n5 IREF.n3 1.33272
R3558 IREF.n73 IREF.n30 1.13717
R3559 IREF.n73 IREF.n72 1.09471
R3560 IREF.n120 IREF.n119 0.438108
R3561 IREF.n97 IREF 0.43525
R3562 IREF.n118 IREF.n117 0.433991
R3563 IREF.n72 IREF.n46 0.374888
R3564 IREF.n30 IREF.n29 0.374529
R3565 IREF.n17 IREF.n16 0.166571
R3566 IREF.n41 IREF.n40 0.166571
R3567 IREF.n65 IREF.n64 0.166571
R3568 IREF.n110 IREF.n103 0.166571
R3569 IREF.n127 IREF.n126 0.166571
R3570 IREF.n91 IREF.n90 0.166571
R3571 IREF.n26 IREF.n25 0.142774
R3572 IREF.n6 IREF.n5 0.139606
R3573 IREF IREF.n133 0.126773
R3574 IREF.n29 IREF.n23 0.114786
R3575 IREF.n9 IREF.n3 0.114786
R3576 IREF.n15 IREF.n10 0.114786
R3577 IREF.n16 IREF.n15 0.114786
R3578 IREF.n17 IREF.n0 0.114786
R3579 IREF.n22 IREF.n0 0.114786
R3580 IREF.n46 IREF.n31 0.114786
R3581 IREF.n41 IREF.n31 0.114786
R3582 IREF.n40 IREF.n39 0.114786
R3583 IREF.n57 IREF.n50 0.114786
R3584 IREF.n63 IREF.n58 0.114786
R3585 IREF.n64 IREF.n63 0.114786
R3586 IREF.n65 IREF.n47 0.114786
R3587 IREF.n71 IREF.n47 0.114786
R3588 IREF.n116 IREF.n103 0.114786
R3589 IREF.n110 IREF.n109 0.114786
R3590 IREF.n109 IREF.n105 0.114786
R3591 IREF.n125 IREF.n101 0.114786
R3592 IREF.n126 IREF.n125 0.114786
R3593 IREF.n127 IREF.n98 0.114786
R3594 IREF.n132 IREF.n98 0.114786
R3595 IREF.n83 IREF.n77 0.114786
R3596 IREF.n89 IREF.n84 0.114786
R3597 IREF.n90 IREF.n89 0.114786
R3598 IREF.n91 IREF.n74 0.114786
R3599 IREF.n96 IREF.n74 0.114786
R3600 IREF.n18 IREF.n2 0.0899231
R3601 IREF.n128 IREF.n100 0.0899231
R3602 IREF.n112 IREF.n111 0.0899231
R3603 IREF.n80 IREF.n79 0.0669267
R3604 IREF.n53 IREF.n52 0.0662833
R3605 IREF.n28 IREF.n24 0.0572308
R3606 IREF.n108 IREF.n107 0.0553077
R3607 IREF.n131 IREF.n99 0.0543462
R3608 IREF.n21 IREF.n1 0.0533846
R3609 IREF.n14 IREF.n11 0.0524231
R3610 IREF.n8 IREF.n4 0.0524231
R3611 IREF.n124 IREF.n121 0.0514615
R3612 IREF.n115 IREF.n102 0.0505
R3613 IREF.n111 IREF.n104 0.0476154
R3614 IREF IREF.n73 0.0475
R3615 IREF.n129 IREF.n128 0.0466538
R3616 IREF.n19 IREF.n18 0.0456923
R3617 IREF.n13 IREF.n2 0.0447308
R3618 IREF.n123 IREF.n100 0.0437692
R3619 IREF.n133 IREF.n97 0.0429567
R3620 IREF.n114 IREF.n112 0.0428077
R3621 IREF.n42 IREF.n33 0.0420179
R3622 IREF.n66 IREF.n49 0.0420179
R3623 IREF.n92 IREF.n76 0.0418701
R3624 IREF.n45 IREF.n32 0.0268393
R3625 IREF.n82 IREF.n78 0.0258559
R3626 IREF.n95 IREF.n75 0.025411
R3627 IREF.n69 IREF.n48 0.0250536
R3628 IREF.n62 IREF.n59 0.0246071
R3629 IREF.n55 IREF.n51 0.0246071
R3630 IREF.n88 IREF.n85 0.0240765
R3631 IREF.n43 IREF.n42 0.0232679
R3632 IREF.n38 IREF.n37 0.0228214
R3633 IREF.n93 IREF.n92 0.0218523
R3634 IREF.n67 IREF.n66 0.0214821
R3635 IREF.n61 IREF.n49 0.0210357
R3636 IREF.n87 IREF.n76 0.0205178
R3637 IREF.n115 IREF.n114 0.0197308
R3638 IREF.n35 IREF.n33 0.01925
R3639 IREF.n124 IREF.n123 0.0187692
R3640 IREF.n14 IREF.n13 0.0178077
R3641 IREF.n6 IREF.n4 0.0178077
R3642 IREF.n19 IREF.n1 0.0168462
R3643 IREF.n129 IREF.n99 0.0158846
R3644 IREF.n108 IREF.n104 0.0149231
R3645 IREF.n26 IREF.n24 0.013
R3646 IREF.n117 IREF.n102 0.0120385
R3647 IREF.n121 IREF.n120 0.0110769
R3648 IREF.n38 IREF.n35 0.0103214
R3649 IREF.n88 IREF.n87 0.00895196
R3650 IREF.n62 IREF.n61 0.00853571
R3651 IREF.n53 IREF.n51 0.00853571
R3652 IREF.n67 IREF.n48 0.00808929
R3653 IREF.n93 IREF.n75 0.00761744
R3654 IREF.n80 IREF.n78 0.0071726
R3655 IREF.n37 IREF.n34 0.00675
R3656 IREF.n43 IREF.n32 0.00630357
R3657 IREF.n56 IREF.n55 0.00496429
R3658 IREF.n70 IREF.n69 0.00451786
R3659 VB1.n174 VB1.t44 233.504
R3660 VB1.n337 VB1.t52 232.321
R3661 VB1.n255 VB1.t40 232.317
R3662 VB1.n337 VB1.t68 231.948
R3663 VB1.n255 VB1.t20 231.946
R3664 VB1.n173 VB1.n171 207.048
R3665 VB1.n175 VB1.n170 205.881
R3666 VB1.n173 VB1.n172 204.861
R3667 VB1.n329 VB1.n327 203.756
R3668 VB1.n335 VB1.n333 203.756
R3669 VB1.n332 VB1.n331 203.756
R3670 VB1.n247 VB1.n245 203.752
R3671 VB1.n253 VB1.n251 203.752
R3672 VB1.n250 VB1.n249 203.752
R3673 VB1.n329 VB1.n328 203.383
R3674 VB1.n335 VB1.n334 203.383
R3675 VB1.n332 VB1.n330 203.383
R3676 VB1.n247 VB1.n246 203.381
R3677 VB1.n253 VB1.n252 203.381
R3678 VB1.n250 VB1.n248 203.381
R3679 VB1.n45 VB1.t242 113.686
R3680 VB1.n113 VB1.t111 113.686
R3681 VB1.n140 VB1.t120 113.686
R3682 VB1.n188 VB1.t171 113.686
R3683 VB1.n215 VB1.t200 113.686
R3684 VB1.n297 VB1.t84 113.686
R3685 VB1.n352 VB1.t201 113.686
R3686 VB1.n453 VB1.t157 113.686
R3687 VB1.n4 VB1.t156 113.686
R3688 VB1.n72 VB1.t191 113.686
R3689 VB1.n379 VB1.t179 113.686
R3690 VB1.n413 VB1.t86 113.686
R3691 VB1.n270 VB1.t245 113.684
R3692 VB1.n35 VB1.t159 113.683
R3693 VB1.n103 VB1.t206 113.683
R3694 VB1.n162 VB1.t219 113.683
R3695 VB1.n178 VB1.t59 113.683
R3696 VB1.n237 VB1.t31 113.683
R3697 VB1.n319 VB1.t37 113.683
R3698 VB1.n342 VB1.t47 113.683
R3699 VB1.n478 VB1.t103 113.683
R3700 VB1.n443 VB1.t226 113.683
R3701 VB1.n26 VB1.t87 113.681
R3702 VB1.n94 VB1.t122 113.681
R3703 VB1.n401 VB1.t229 113.681
R3704 VB1.n495 VB1.t175 113.681
R3705 VB1.n435 VB1.t150 113.681
R3706 VB1.n260 VB1.t25 113.681
R3707 VB1.n35 VB1.t161 113.68
R3708 VB1.n103 VB1.t209 113.68
R3709 VB1.n162 VB1.t221 113.68
R3710 VB1.n178 VB1.t109 113.68
R3711 VB1.n237 VB1.t128 113.68
R3712 VB1.n319 VB1.t188 113.68
R3713 VB1.n342 VB1.t115 113.68
R3714 VB1.n478 VB1.t106 113.68
R3715 VB1.n443 VB1.t170 113.68
R3716 VB1.n26 VB1.t92 113.677
R3717 VB1.n94 VB1.t127 113.677
R3718 VB1.n401 VB1.t93 113.677
R3719 VB1.n495 VB1.t134 113.677
R3720 VB1.n435 VB1.t102 113.677
R3721 VB1.n260 VB1.t164 113.677
R3722 VB1.n45 VB1.t233 113.675
R3723 VB1.n113 VB1.t94 113.675
R3724 VB1.n140 VB1.t112 113.675
R3725 VB1.n188 VB1.t41 113.675
R3726 VB1.n215 VB1.t9 113.675
R3727 VB1.n297 VB1.t65 113.675
R3728 VB1.n352 VB1.t55 113.675
R3729 VB1.n453 VB1.t85 113.675
R3730 VB1.n4 VB1.t152 113.674
R3731 VB1.n72 VB1.t177 113.674
R3732 VB1.n379 VB1.t82 113.674
R3733 VB1.n413 VB1.t183 113.674
R3734 VB1.n270 VB1.t29 113.674
R3735 VB1.n39 VB1.t80 113.624
R3736 VB1.n62 VB1.t81 113.624
R3737 VB1.n57 VB1.t139 113.624
R3738 VB1.n52 VB1.t135 113.624
R3739 VB1.n47 VB1.t187 113.624
R3740 VB1.n107 VB1.t130 113.624
R3741 VB1.n130 VB1.t129 113.624
R3742 VB1.n125 VB1.t174 113.624
R3743 VB1.n120 VB1.t160 113.624
R3744 VB1.n115 VB1.t230 113.624
R3745 VB1.n166 VB1.t141 113.624
R3746 VB1.n157 VB1.t140 113.624
R3747 VB1.n152 VB1.t186 113.624
R3748 VB1.n147 VB1.t176 113.624
R3749 VB1.n142 VB1.t244 113.624
R3750 VB1.n182 VB1.t196 113.624
R3751 VB1.n205 VB1.t195 113.624
R3752 VB1.n200 VB1.t13 113.624
R3753 VB1.n195 VB1.t241 113.624
R3754 VB1.n190 VB1.t61 113.624
R3755 VB1.n241 VB1.t218 113.624
R3756 VB1.n232 VB1.t217 113.624
R3757 VB1.n227 VB1.t69 113.624
R3758 VB1.n222 VB1.t79 113.624
R3759 VB1.n217 VB1.t11 113.624
R3760 VB1.n323 VB1.t114 113.624
R3761 VB1.n314 VB1.t113 113.624
R3762 VB1.n309 VB1.t15 113.624
R3763 VB1.n304 VB1.t151 113.624
R3764 VB1.n299 VB1.t21 113.624
R3765 VB1.n346 VB1.t248 113.624
R3766 VB1.n369 VB1.t185 113.624
R3767 VB1.n364 VB1.t45 113.624
R3768 VB1.n359 VB1.t124 113.624
R3769 VB1.n354 VB1.t33 113.624
R3770 VB1.n482 VB1.t193 113.624
R3771 VB1.n553 VB1.t192 113.624
R3772 VB1.n548 VB1.t246 113.624
R3773 VB1.n543 VB1.t240 113.624
R3774 VB1.n538 VB1.t126 113.624
R3775 VB1.n533 VB1.t165 113.624
R3776 VB1.n447 VB1.t249 113.624
R3777 VB1.n470 VB1.t99 113.624
R3778 VB1.n465 VB1.t158 113.624
R3779 VB1.n460 VB1.t95 113.624
R3780 VB1.n455 VB1.t98 113.624
R3781 VB1.n30 VB1.t180 113.624
R3782 VB1.n21 VB1.t181 113.624
R3783 VB1.n16 VB1.t239 113.624
R3784 VB1.n11 VB1.t231 113.624
R3785 VB1.n6 VB1.t117 113.624
R3786 VB1.n98 VB1.t213 113.624
R3787 VB1.n89 VB1.t212 113.624
R3788 VB1.n84 VB1.t91 113.624
R3789 VB1.n79 VB1.t76 113.624
R3790 VB1.n74 VB1.t144 113.624
R3791 VB1.n405 VB1.t238 113.624
R3792 VB1.n396 VB1.t163 113.624
R3793 VB1.n391 VB1.t178 113.624
R3794 VB1.n386 VB1.t108 113.624
R3795 VB1.n381 VB1.t168 113.624
R3796 VB1.n505 VB1.t225 113.624
R3797 VB1.n510 VB1.t123 113.624
R3798 VB1.n515 VB1.t223 113.624
R3799 VB1.n520 VB1.t224 113.624
R3800 VB1.n525 VB1.t121 113.624
R3801 VB1.n499 VB1.t205 113.624
R3802 VB1.n439 VB1.t172 113.624
R3803 VB1.n430 VB1.t198 113.624
R3804 VB1.n425 VB1.t88 113.624
R3805 VB1.n420 VB1.t190 113.624
R3806 VB1.n415 VB1.t194 113.624
R3807 VB1.n264 VB1.t90 113.623
R3808 VB1.n287 VB1.t89 113.623
R3809 VB1.n282 VB1.t57 113.623
R3810 VB1.n277 VB1.t136 113.623
R3811 VB1.n272 VB1.t35 113.623
R3812 VB1.n37 VB1.t154 113.617
R3813 VB1.n64 VB1.t222 113.617
R3814 VB1.n59 VB1.t101 113.617
R3815 VB1.n54 VB1.t137 113.617
R3816 VB1.n49 VB1.t189 113.617
R3817 VB1.n105 VB1.t202 113.617
R3818 VB1.n132 VB1.t77 113.617
R3819 VB1.n127 VB1.t138 113.617
R3820 VB1.n122 VB1.t169 113.617
R3821 VB1.n117 VB1.t235 113.617
R3822 VB1.n164 VB1.t211 113.617
R3823 VB1.n159 VB1.t104 113.617
R3824 VB1.n154 VB1.t149 113.617
R3825 VB1.n149 VB1.t182 113.617
R3826 VB1.n144 VB1.t247 113.617
R3827 VB1.n180 VB1.t17 113.617
R3828 VB1.n207 VB1.t43 113.617
R3829 VB1.n202 VB1.t208 113.617
R3830 VB1.n197 VB1.t23 113.617
R3831 VB1.n192 VB1.t133 113.617
R3832 VB1.n239 VB1.t63 113.617
R3833 VB1.n234 VB1.t39 113.617
R3834 VB1.n229 VB1.t228 113.617
R3835 VB1.n224 VB1.t5 113.617
R3836 VB1.n219 VB1.t148 113.617
R3837 VB1.n321 VB1.t49 113.617
R3838 VB1.n316 VB1.t51 113.617
R3839 VB1.n311 VB1.t125 113.617
R3840 VB1.n306 VB1.t53 113.617
R3841 VB1.n301 VB1.t214 113.617
R3842 VB1.n344 VB1.t27 113.617
R3843 VB1.n371 VB1.t67 113.617
R3844 VB1.n366 VB1.t116 113.617
R3845 VB1.n361 VB1.t73 113.617
R3846 VB1.n356 VB1.t232 113.617
R3847 VB1.n480 VB1.t96 113.617
R3848 VB1.n555 VB1.t153 113.617
R3849 VB1.n550 VB1.t207 113.617
R3850 VB1.n545 VB1.t243 113.617
R3851 VB1.n540 VB1.t131 113.617
R3852 VB1.n535 VB1.t155 113.617
R3853 VB1.n445 VB1.t107 113.617
R3854 VB1.n472 VB1.t110 113.617
R3855 VB1.n467 VB1.t167 113.617
R3856 VB1.n462 VB1.t216 113.617
R3857 VB1.n457 VB1.t220 113.617
R3858 VB1.n28 VB1.t78 113.615
R3859 VB1.n23 VB1.t146 113.615
R3860 VB1.n18 VB1.t197 113.615
R3861 VB1.n13 VB1.t236 113.615
R3862 VB1.n8 VB1.t119 113.615
R3863 VB1.n96 VB1.t118 113.615
R3864 VB1.n91 VB1.t173 113.615
R3865 VB1.n86 VB1.t227 113.615
R3866 VB1.n81 VB1.t83 113.615
R3867 VB1.n76 VB1.t147 113.615
R3868 VB1.n403 VB1.t184 113.615
R3869 VB1.n398 VB1.t75 113.615
R3870 VB1.n393 VB1.t97 113.615
R3871 VB1.n388 VB1.t145 113.615
R3872 VB1.n383 VB1.t210 113.615
R3873 VB1.n503 VB1.t237 113.615
R3874 VB1.n508 VB1.t132 113.615
R3875 VB1.n513 VB1.t162 113.615
R3876 VB1.n518 VB1.t166 113.615
R3877 VB1.n523 VB1.t215 113.615
R3878 VB1.n497 VB1.t234 113.615
R3879 VB1.n437 VB1.t203 113.615
R3880 VB1.n432 VB1.t204 113.615
R3881 VB1.n427 VB1.t100 113.615
R3882 VB1.n422 VB1.t142 113.615
R3883 VB1.n417 VB1.t143 113.615
R3884 VB1.n262 VB1.t7 113.615
R3885 VB1.n289 VB1.t19 113.615
R3886 VB1.n284 VB1.t105 113.615
R3887 VB1.n279 VB1.t71 113.615
R3888 VB1.n274 VB1.t199 113.615
R3889 VB1.n529 VB1.t3 92.0321
R3890 VB1.n527 VB1.t1 91.9752
R3891 VB1.n528 VB1.t0 91.5354
R3892 VB1.n529 VB1.t2 89.497
R3893 VB1.n527 VB1.t4 88.9416
R3894 VB1.n170 VB1.t18 28.5655
R3895 VB1.n170 VB1.t60 28.5655
R3896 VB1.n172 VB1.t24 28.5655
R3897 VB1.n172 VB1.t14 28.5655
R3898 VB1.n171 VB1.t42 28.5655
R3899 VB1.n171 VB1.t62 28.5655
R3900 VB1.n246 VB1.t8 28.5655
R3901 VB1.n246 VB1.t26 28.5655
R3902 VB1.n245 VB1.t64 28.5655
R3903 VB1.n245 VB1.t32 28.5655
R3904 VB1.n252 VB1.t72 28.5655
R3905 VB1.n252 VB1.t58 28.5655
R3906 VB1.n251 VB1.t6 28.5655
R3907 VB1.n251 VB1.t70 28.5655
R3908 VB1.n249 VB1.t10 28.5655
R3909 VB1.n249 VB1.t12 28.5655
R3910 VB1.n248 VB1.t30 28.5655
R3911 VB1.n248 VB1.t36 28.5655
R3912 VB1.n328 VB1.t28 28.5655
R3913 VB1.n328 VB1.t48 28.5655
R3914 VB1.n327 VB1.t50 28.5655
R3915 VB1.n327 VB1.t38 28.5655
R3916 VB1.n334 VB1.t74 28.5655
R3917 VB1.n334 VB1.t46 28.5655
R3918 VB1.n333 VB1.t54 28.5655
R3919 VB1.n333 VB1.t16 28.5655
R3920 VB1.n331 VB1.t66 28.5655
R3921 VB1.n331 VB1.t22 28.5655
R3922 VB1.n330 VB1.t56 28.5655
R3923 VB1.n330 VB1.t34 28.5655
R3924 VB1.n28 VB1.n27 4.5005
R3925 VB1.n29 VB1.n25 4.5005
R3926 VB1.n31 VB1.n30 4.5005
R3927 VB1.n9 VB1.n8 4.5005
R3928 VB1.n7 VB1.n3 4.5005
R3929 VB1.n6 VB1.n5 4.5005
R3930 VB1.n14 VB1.n13 4.5005
R3931 VB1.n12 VB1.n2 4.5005
R3932 VB1.n11 VB1.n10 4.5005
R3933 VB1.n19 VB1.n18 4.5005
R3934 VB1.n17 VB1.n1 4.5005
R3935 VB1.n16 VB1.n15 4.5005
R3936 VB1.n24 VB1.n23 4.5005
R3937 VB1.n22 VB1.n0 4.5005
R3938 VB1.n21 VB1.n20 4.5005
R3939 VB1.n37 VB1.n36 4.5005
R3940 VB1.n38 VB1.n34 4.5005
R3941 VB1.n40 VB1.n39 4.5005
R3942 VB1.n50 VB1.n49 4.5005
R3943 VB1.n48 VB1.n44 4.5005
R3944 VB1.n47 VB1.n46 4.5005
R3945 VB1.n55 VB1.n54 4.5005
R3946 VB1.n53 VB1.n43 4.5005
R3947 VB1.n52 VB1.n51 4.5005
R3948 VB1.n60 VB1.n59 4.5005
R3949 VB1.n58 VB1.n42 4.5005
R3950 VB1.n57 VB1.n56 4.5005
R3951 VB1.n65 VB1.n64 4.5005
R3952 VB1.n63 VB1.n41 4.5005
R3953 VB1.n62 VB1.n61 4.5005
R3954 VB1.n96 VB1.n95 4.5005
R3955 VB1.n97 VB1.n93 4.5005
R3956 VB1.n99 VB1.n98 4.5005
R3957 VB1.n77 VB1.n76 4.5005
R3958 VB1.n75 VB1.n71 4.5005
R3959 VB1.n74 VB1.n73 4.5005
R3960 VB1.n82 VB1.n81 4.5005
R3961 VB1.n80 VB1.n70 4.5005
R3962 VB1.n79 VB1.n78 4.5005
R3963 VB1.n87 VB1.n86 4.5005
R3964 VB1.n85 VB1.n69 4.5005
R3965 VB1.n84 VB1.n83 4.5005
R3966 VB1.n92 VB1.n91 4.5005
R3967 VB1.n90 VB1.n68 4.5005
R3968 VB1.n89 VB1.n88 4.5005
R3969 VB1.n105 VB1.n104 4.5005
R3970 VB1.n106 VB1.n102 4.5005
R3971 VB1.n108 VB1.n107 4.5005
R3972 VB1.n118 VB1.n117 4.5005
R3973 VB1.n116 VB1.n112 4.5005
R3974 VB1.n115 VB1.n114 4.5005
R3975 VB1.n123 VB1.n122 4.5005
R3976 VB1.n121 VB1.n111 4.5005
R3977 VB1.n120 VB1.n119 4.5005
R3978 VB1.n128 VB1.n127 4.5005
R3979 VB1.n126 VB1.n110 4.5005
R3980 VB1.n125 VB1.n124 4.5005
R3981 VB1.n133 VB1.n132 4.5005
R3982 VB1.n131 VB1.n109 4.5005
R3983 VB1.n130 VB1.n129 4.5005
R3984 VB1.n164 VB1.n163 4.5005
R3985 VB1.n165 VB1.n161 4.5005
R3986 VB1.n167 VB1.n166 4.5005
R3987 VB1.n145 VB1.n144 4.5005
R3988 VB1.n143 VB1.n139 4.5005
R3989 VB1.n142 VB1.n141 4.5005
R3990 VB1.n150 VB1.n149 4.5005
R3991 VB1.n148 VB1.n138 4.5005
R3992 VB1.n147 VB1.n146 4.5005
R3993 VB1.n155 VB1.n154 4.5005
R3994 VB1.n153 VB1.n137 4.5005
R3995 VB1.n152 VB1.n151 4.5005
R3996 VB1.n160 VB1.n159 4.5005
R3997 VB1.n158 VB1.n136 4.5005
R3998 VB1.n157 VB1.n156 4.5005
R3999 VB1.n180 VB1.n179 4.5005
R4000 VB1.n181 VB1.n177 4.5005
R4001 VB1.n183 VB1.n182 4.5005
R4002 VB1.n193 VB1.n192 4.5005
R4003 VB1.n191 VB1.n187 4.5005
R4004 VB1.n190 VB1.n189 4.5005
R4005 VB1.n198 VB1.n197 4.5005
R4006 VB1.n196 VB1.n186 4.5005
R4007 VB1.n195 VB1.n194 4.5005
R4008 VB1.n203 VB1.n202 4.5005
R4009 VB1.n201 VB1.n185 4.5005
R4010 VB1.n200 VB1.n199 4.5005
R4011 VB1.n208 VB1.n207 4.5005
R4012 VB1.n206 VB1.n184 4.5005
R4013 VB1.n205 VB1.n204 4.5005
R4014 VB1.n239 VB1.n238 4.5005
R4015 VB1.n240 VB1.n236 4.5005
R4016 VB1.n242 VB1.n241 4.5005
R4017 VB1.n220 VB1.n219 4.5005
R4018 VB1.n218 VB1.n214 4.5005
R4019 VB1.n217 VB1.n216 4.5005
R4020 VB1.n225 VB1.n224 4.5005
R4021 VB1.n223 VB1.n213 4.5005
R4022 VB1.n222 VB1.n221 4.5005
R4023 VB1.n230 VB1.n229 4.5005
R4024 VB1.n228 VB1.n212 4.5005
R4025 VB1.n227 VB1.n226 4.5005
R4026 VB1.n235 VB1.n234 4.5005
R4027 VB1.n233 VB1.n211 4.5005
R4028 VB1.n232 VB1.n231 4.5005
R4029 VB1.n262 VB1.n261 4.5005
R4030 VB1.n263 VB1.n259 4.5005
R4031 VB1.n265 VB1.n264 4.5005
R4032 VB1.n275 VB1.n274 4.5005
R4033 VB1.n273 VB1.n269 4.5005
R4034 VB1.n272 VB1.n271 4.5005
R4035 VB1.n280 VB1.n279 4.5005
R4036 VB1.n278 VB1.n268 4.5005
R4037 VB1.n277 VB1.n276 4.5005
R4038 VB1.n285 VB1.n284 4.5005
R4039 VB1.n283 VB1.n267 4.5005
R4040 VB1.n282 VB1.n281 4.5005
R4041 VB1.n290 VB1.n289 4.5005
R4042 VB1.n288 VB1.n266 4.5005
R4043 VB1.n287 VB1.n286 4.5005
R4044 VB1.n321 VB1.n320 4.5005
R4045 VB1.n322 VB1.n318 4.5005
R4046 VB1.n324 VB1.n323 4.5005
R4047 VB1.n302 VB1.n301 4.5005
R4048 VB1.n300 VB1.n296 4.5005
R4049 VB1.n299 VB1.n298 4.5005
R4050 VB1.n307 VB1.n306 4.5005
R4051 VB1.n305 VB1.n295 4.5005
R4052 VB1.n304 VB1.n303 4.5005
R4053 VB1.n312 VB1.n311 4.5005
R4054 VB1.n310 VB1.n294 4.5005
R4055 VB1.n309 VB1.n308 4.5005
R4056 VB1.n317 VB1.n316 4.5005
R4057 VB1.n315 VB1.n293 4.5005
R4058 VB1.n314 VB1.n313 4.5005
R4059 VB1.n344 VB1.n343 4.5005
R4060 VB1.n345 VB1.n341 4.5005
R4061 VB1.n347 VB1.n346 4.5005
R4062 VB1.n357 VB1.n356 4.5005
R4063 VB1.n355 VB1.n351 4.5005
R4064 VB1.n354 VB1.n353 4.5005
R4065 VB1.n362 VB1.n361 4.5005
R4066 VB1.n360 VB1.n350 4.5005
R4067 VB1.n359 VB1.n358 4.5005
R4068 VB1.n367 VB1.n366 4.5005
R4069 VB1.n365 VB1.n349 4.5005
R4070 VB1.n364 VB1.n363 4.5005
R4071 VB1.n372 VB1.n371 4.5005
R4072 VB1.n370 VB1.n348 4.5005
R4073 VB1.n369 VB1.n368 4.5005
R4074 VB1.n403 VB1.n402 4.5005
R4075 VB1.n404 VB1.n400 4.5005
R4076 VB1.n406 VB1.n405 4.5005
R4077 VB1.n384 VB1.n383 4.5005
R4078 VB1.n382 VB1.n378 4.5005
R4079 VB1.n381 VB1.n380 4.5005
R4080 VB1.n389 VB1.n388 4.5005
R4081 VB1.n387 VB1.n377 4.5005
R4082 VB1.n386 VB1.n385 4.5005
R4083 VB1.n394 VB1.n393 4.5005
R4084 VB1.n392 VB1.n376 4.5005
R4085 VB1.n391 VB1.n390 4.5005
R4086 VB1.n399 VB1.n398 4.5005
R4087 VB1.n397 VB1.n375 4.5005
R4088 VB1.n396 VB1.n395 4.5005
R4089 VB1.n480 VB1.n479 4.5005
R4090 VB1.n481 VB1.n477 4.5005
R4091 VB1.n483 VB1.n482 4.5005
R4092 VB1.n497 VB1.n496 4.5005
R4093 VB1.n498 VB1.n494 4.5005
R4094 VB1.n500 VB1.n499 4.5005
R4095 VB1.n523 VB1.n522 4.5005
R4096 VB1.n524 VB1.n489 4.5005
R4097 VB1.n526 VB1.n525 4.5005
R4098 VB1.n518 VB1.n517 4.5005
R4099 VB1.n519 VB1.n490 4.5005
R4100 VB1.n521 VB1.n520 4.5005
R4101 VB1.n513 VB1.n512 4.5005
R4102 VB1.n514 VB1.n491 4.5005
R4103 VB1.n516 VB1.n515 4.5005
R4104 VB1.n508 VB1.n507 4.5005
R4105 VB1.n509 VB1.n492 4.5005
R4106 VB1.n511 VB1.n510 4.5005
R4107 VB1.n503 VB1.n502 4.5005
R4108 VB1.n504 VB1.n493 4.5005
R4109 VB1.n506 VB1.n505 4.5005
R4110 VB1.n536 VB1.n535 4.5005
R4111 VB1.n534 VB1.n488 4.5005
R4112 VB1.n533 VB1.n532 4.5005
R4113 VB1.n541 VB1.n540 4.5005
R4114 VB1.n539 VB1.n487 4.5005
R4115 VB1.n538 VB1.n537 4.5005
R4116 VB1.n546 VB1.n545 4.5005
R4117 VB1.n544 VB1.n486 4.5005
R4118 VB1.n543 VB1.n542 4.5005
R4119 VB1.n551 VB1.n550 4.5005
R4120 VB1.n549 VB1.n485 4.5005
R4121 VB1.n548 VB1.n547 4.5005
R4122 VB1.n556 VB1.n555 4.5005
R4123 VB1.n554 VB1.n484 4.5005
R4124 VB1.n553 VB1.n552 4.5005
R4125 VB1.n445 VB1.n444 4.5005
R4126 VB1.n446 VB1.n442 4.5005
R4127 VB1.n448 VB1.n447 4.5005
R4128 VB1.n458 VB1.n457 4.5005
R4129 VB1.n456 VB1.n452 4.5005
R4130 VB1.n455 VB1.n454 4.5005
R4131 VB1.n463 VB1.n462 4.5005
R4132 VB1.n461 VB1.n451 4.5005
R4133 VB1.n460 VB1.n459 4.5005
R4134 VB1.n468 VB1.n467 4.5005
R4135 VB1.n466 VB1.n450 4.5005
R4136 VB1.n465 VB1.n464 4.5005
R4137 VB1.n473 VB1.n472 4.5005
R4138 VB1.n471 VB1.n449 4.5005
R4139 VB1.n470 VB1.n469 4.5005
R4140 VB1.n437 VB1.n436 4.5005
R4141 VB1.n438 VB1.n434 4.5005
R4142 VB1.n440 VB1.n439 4.5005
R4143 VB1.n418 VB1.n417 4.5005
R4144 VB1.n416 VB1.n412 4.5005
R4145 VB1.n415 VB1.n414 4.5005
R4146 VB1.n423 VB1.n422 4.5005
R4147 VB1.n421 VB1.n411 4.5005
R4148 VB1.n420 VB1.n419 4.5005
R4149 VB1.n428 VB1.n427 4.5005
R4150 VB1.n426 VB1.n410 4.5005
R4151 VB1.n425 VB1.n424 4.5005
R4152 VB1.n433 VB1.n432 4.5005
R4153 VB1.n431 VB1.n409 4.5005
R4154 VB1.n430 VB1.n429 4.5005
R4155 VB1.n531 VB1.n526 3.81657
R4156 VB1.n532 VB1.n531 3.81657
R4157 VB1.n254 VB1.n250 3.66453
R4158 VB1.n336 VB1.n332 3.66453
R4159 VB1.n257 VB1.n247 2.49802
R4160 VB1.n339 VB1.n329 2.49802
R4161 VB1.n271 VB1.n270 2.22976
R4162 VB1.n261 VB1.n260 2.22976
R4163 VB1.n5 VB1.n4 2.22967
R4164 VB1.n73 VB1.n72 2.22967
R4165 VB1.n380 VB1.n379 2.22967
R4166 VB1.n414 VB1.n413 2.22967
R4167 VB1.n27 VB1.n26 2.22967
R4168 VB1.n95 VB1.n94 2.22967
R4169 VB1.n402 VB1.n401 2.22967
R4170 VB1.n496 VB1.n495 2.22967
R4171 VB1.n436 VB1.n435 2.22967
R4172 VB1.n36 VB1.n35 2.22939
R4173 VB1.n46 VB1.n45 2.22939
R4174 VB1.n104 VB1.n103 2.22939
R4175 VB1.n114 VB1.n113 2.22939
R4176 VB1.n163 VB1.n162 2.22939
R4177 VB1.n141 VB1.n140 2.22939
R4178 VB1.n179 VB1.n178 2.22939
R4179 VB1.n189 VB1.n188 2.22939
R4180 VB1.n238 VB1.n237 2.22939
R4181 VB1.n216 VB1.n215 2.22939
R4182 VB1.n320 VB1.n319 2.22939
R4183 VB1.n298 VB1.n297 2.22939
R4184 VB1.n343 VB1.n342 2.22939
R4185 VB1.n353 VB1.n352 2.22939
R4186 VB1.n479 VB1.n478 2.22939
R4187 VB1.n444 VB1.n443 2.22939
R4188 VB1.n454 VB1.n453 2.22939
R4189 VB1.n531 VB1.n530 2.04075
R4190 VB1.n174 VB1.n173 1.68288
R4191 VB1.n338 VB1.n336 1.68288
R4192 VB1.n256 VB1.n254 1.6808
R4193 VB1.n256 VB1.n255 1.55537
R4194 VB1.n338 VB1.n337 1.55537
R4195 VB1.n254 VB1.n253 1.47765
R4196 VB1.n336 VB1.n335 1.47765
R4197 VB1 VB1.n528 1.30934
R4198 VB1.n475 VB1.n441 1.12134
R4199 VB1.n530 VB1.n529 1.0963
R4200 VB1.n475 VB1.n474 1.09471
R4201 VB1.n558 VB1.n557 1.09471
R4202 VB1.n501 VB1.n476 1.09471
R4203 VB1.n408 VB1.n407 1.09471
R4204 VB1.n374 VB1.n373 1.09471
R4205 VB1.n326 VB1.n325 1.09471
R4206 VB1.n292 VB1.n291 1.09471
R4207 VB1.n244 VB1.n243 1.09471
R4208 VB1.n210 VB1.n209 1.09471
R4209 VB1.n169 VB1.n168 1.09471
R4210 VB1.n135 VB1.n134 1.09471
R4211 VB1.n101 VB1.n100 1.09471
R4212 VB1.n67 VB1.n66 1.09471
R4213 VB1.n33 VB1.n32 1.09471
R4214 VB1.n340 VB1.n339 1.09471
R4215 VB1.n258 VB1.n257 1.09471
R4216 VB1.n176 VB1.n175 1.09471
R4217 VB1.n10 VB1.n9 1.03979
R4218 VB1.n51 VB1.n50 1.03979
R4219 VB1.n78 VB1.n77 1.03979
R4220 VB1.n119 VB1.n118 1.03979
R4221 VB1.n146 VB1.n145 1.03979
R4222 VB1.n194 VB1.n193 1.03979
R4223 VB1.n221 VB1.n220 1.03979
R4224 VB1.n276 VB1.n275 1.03979
R4225 VB1.n303 VB1.n302 1.03979
R4226 VB1.n358 VB1.n357 1.03979
R4227 VB1.n385 VB1.n384 1.03979
R4228 VB1.n517 VB1.n516 1.03979
R4229 VB1.n542 VB1.n541 1.03979
R4230 VB1.n459 VB1.n458 1.03979
R4231 VB1.n419 VB1.n418 1.03979
R4232 VB1.n15 VB1.n14 0.693357
R4233 VB1.n20 VB1.n19 0.693357
R4234 VB1.n56 VB1.n55 0.693357
R4235 VB1.n61 VB1.n60 0.693357
R4236 VB1.n83 VB1.n82 0.693357
R4237 VB1.n88 VB1.n87 0.693357
R4238 VB1.n124 VB1.n123 0.693357
R4239 VB1.n129 VB1.n128 0.693357
R4240 VB1.n151 VB1.n150 0.693357
R4241 VB1.n156 VB1.n155 0.693357
R4242 VB1.n199 VB1.n198 0.693357
R4243 VB1.n204 VB1.n203 0.693357
R4244 VB1.n226 VB1.n225 0.693357
R4245 VB1.n231 VB1.n230 0.693357
R4246 VB1.n281 VB1.n280 0.693357
R4247 VB1.n286 VB1.n285 0.693357
R4248 VB1.n308 VB1.n307 0.693357
R4249 VB1.n313 VB1.n312 0.693357
R4250 VB1.n363 VB1.n362 0.693357
R4251 VB1.n368 VB1.n367 0.693357
R4252 VB1.n390 VB1.n389 0.693357
R4253 VB1.n395 VB1.n394 0.693357
R4254 VB1.n522 VB1.n521 0.693357
R4255 VB1.n512 VB1.n511 0.693357
R4256 VB1.n507 VB1.n506 0.693357
R4257 VB1.n537 VB1.n536 0.693357
R4258 VB1.n547 VB1.n546 0.693357
R4259 VB1.n552 VB1.n551 0.693357
R4260 VB1.n464 VB1.n463 0.693357
R4261 VB1.n469 VB1.n468 0.693357
R4262 VB1.n424 VB1.n423 0.693357
R4263 VB1.n429 VB1.n428 0.693357
R4264 VB1.n66 VB1.n40 0.451674
R4265 VB1.n134 VB1.n108 0.451674
R4266 VB1.n209 VB1.n183 0.451674
R4267 VB1.n291 VB1.n265 0.451674
R4268 VB1.n373 VB1.n347 0.451674
R4269 VB1.n557 VB1.n483 0.451674
R4270 VB1.n474 VB1.n448 0.451674
R4271 VB1.n32 VB1.n31 0.451315
R4272 VB1.n100 VB1.n99 0.451315
R4273 VB1.n168 VB1.n167 0.451315
R4274 VB1.n243 VB1.n242 0.451315
R4275 VB1.n325 VB1.n324 0.451315
R4276 VB1.n407 VB1.n406 0.451315
R4277 VB1.n501 VB1.n500 0.451315
R4278 VB1.n441 VB1.n440 0.451315
R4279 VB1.n502 VB1.n501 0.424531
R4280 VB1.n32 VB1.n24 0.424531
R4281 VB1.n100 VB1.n92 0.424531
R4282 VB1.n168 VB1.n160 0.424531
R4283 VB1.n243 VB1.n235 0.424531
R4284 VB1.n325 VB1.n317 0.424531
R4285 VB1.n407 VB1.n399 0.424531
R4286 VB1.n441 VB1.n433 0.424531
R4287 VB1.n66 VB1.n65 0.424172
R4288 VB1.n134 VB1.n133 0.424172
R4289 VB1.n209 VB1.n208 0.424172
R4290 VB1.n291 VB1.n290 0.424172
R4291 VB1.n373 VB1.n372 0.424172
R4292 VB1.n557 VB1.n556 0.424172
R4293 VB1.n474 VB1.n473 0.424172
R4294 VB1.n528 VB1.n527 0.289473
R4295 VB1.n175 VB1.n174 0.239726
R4296 VB1.n257 VB1.n256 0.239726
R4297 VB1.n339 VB1.n338 0.239726
R4298 VB1.n530 VB1 0.223907
R4299 VB1.n67 VB1.n33 0.209493
R4300 VB1.n135 VB1.n101 0.209493
R4301 VB1.n476 VB1.n475 0.209493
R4302 VB1 VB1.n408 0.133823
R4303 VB1.n176 VB1.n169 0.128653
R4304 VB1.n31 VB1.n25 0.114786
R4305 VB1.n27 VB1.n25 0.114786
R4306 VB1.n5 VB1.n3 0.114786
R4307 VB1.n9 VB1.n3 0.114786
R4308 VB1.n10 VB1.n2 0.114786
R4309 VB1.n14 VB1.n2 0.114786
R4310 VB1.n15 VB1.n1 0.114786
R4311 VB1.n19 VB1.n1 0.114786
R4312 VB1.n20 VB1.n0 0.114786
R4313 VB1.n24 VB1.n0 0.114786
R4314 VB1.n40 VB1.n34 0.114786
R4315 VB1.n36 VB1.n34 0.114786
R4316 VB1.n46 VB1.n44 0.114786
R4317 VB1.n50 VB1.n44 0.114786
R4318 VB1.n51 VB1.n43 0.114786
R4319 VB1.n55 VB1.n43 0.114786
R4320 VB1.n56 VB1.n42 0.114786
R4321 VB1.n60 VB1.n42 0.114786
R4322 VB1.n61 VB1.n41 0.114786
R4323 VB1.n65 VB1.n41 0.114786
R4324 VB1.n99 VB1.n93 0.114786
R4325 VB1.n95 VB1.n93 0.114786
R4326 VB1.n73 VB1.n71 0.114786
R4327 VB1.n77 VB1.n71 0.114786
R4328 VB1.n78 VB1.n70 0.114786
R4329 VB1.n82 VB1.n70 0.114786
R4330 VB1.n83 VB1.n69 0.114786
R4331 VB1.n87 VB1.n69 0.114786
R4332 VB1.n88 VB1.n68 0.114786
R4333 VB1.n92 VB1.n68 0.114786
R4334 VB1.n108 VB1.n102 0.114786
R4335 VB1.n104 VB1.n102 0.114786
R4336 VB1.n114 VB1.n112 0.114786
R4337 VB1.n118 VB1.n112 0.114786
R4338 VB1.n119 VB1.n111 0.114786
R4339 VB1.n123 VB1.n111 0.114786
R4340 VB1.n124 VB1.n110 0.114786
R4341 VB1.n128 VB1.n110 0.114786
R4342 VB1.n129 VB1.n109 0.114786
R4343 VB1.n133 VB1.n109 0.114786
R4344 VB1.n167 VB1.n161 0.114786
R4345 VB1.n163 VB1.n161 0.114786
R4346 VB1.n141 VB1.n139 0.114786
R4347 VB1.n145 VB1.n139 0.114786
R4348 VB1.n146 VB1.n138 0.114786
R4349 VB1.n150 VB1.n138 0.114786
R4350 VB1.n151 VB1.n137 0.114786
R4351 VB1.n155 VB1.n137 0.114786
R4352 VB1.n156 VB1.n136 0.114786
R4353 VB1.n160 VB1.n136 0.114786
R4354 VB1.n183 VB1.n177 0.114786
R4355 VB1.n179 VB1.n177 0.114786
R4356 VB1.n189 VB1.n187 0.114786
R4357 VB1.n193 VB1.n187 0.114786
R4358 VB1.n194 VB1.n186 0.114786
R4359 VB1.n198 VB1.n186 0.114786
R4360 VB1.n199 VB1.n185 0.114786
R4361 VB1.n203 VB1.n185 0.114786
R4362 VB1.n204 VB1.n184 0.114786
R4363 VB1.n208 VB1.n184 0.114786
R4364 VB1.n242 VB1.n236 0.114786
R4365 VB1.n238 VB1.n236 0.114786
R4366 VB1.n216 VB1.n214 0.114786
R4367 VB1.n220 VB1.n214 0.114786
R4368 VB1.n221 VB1.n213 0.114786
R4369 VB1.n225 VB1.n213 0.114786
R4370 VB1.n226 VB1.n212 0.114786
R4371 VB1.n230 VB1.n212 0.114786
R4372 VB1.n231 VB1.n211 0.114786
R4373 VB1.n235 VB1.n211 0.114786
R4374 VB1.n265 VB1.n259 0.114786
R4375 VB1.n261 VB1.n259 0.114786
R4376 VB1.n271 VB1.n269 0.114786
R4377 VB1.n275 VB1.n269 0.114786
R4378 VB1.n276 VB1.n268 0.114786
R4379 VB1.n280 VB1.n268 0.114786
R4380 VB1.n281 VB1.n267 0.114786
R4381 VB1.n285 VB1.n267 0.114786
R4382 VB1.n286 VB1.n266 0.114786
R4383 VB1.n290 VB1.n266 0.114786
R4384 VB1.n324 VB1.n318 0.114786
R4385 VB1.n320 VB1.n318 0.114786
R4386 VB1.n298 VB1.n296 0.114786
R4387 VB1.n302 VB1.n296 0.114786
R4388 VB1.n303 VB1.n295 0.114786
R4389 VB1.n307 VB1.n295 0.114786
R4390 VB1.n308 VB1.n294 0.114786
R4391 VB1.n312 VB1.n294 0.114786
R4392 VB1.n313 VB1.n293 0.114786
R4393 VB1.n317 VB1.n293 0.114786
R4394 VB1.n347 VB1.n341 0.114786
R4395 VB1.n343 VB1.n341 0.114786
R4396 VB1.n353 VB1.n351 0.114786
R4397 VB1.n357 VB1.n351 0.114786
R4398 VB1.n358 VB1.n350 0.114786
R4399 VB1.n362 VB1.n350 0.114786
R4400 VB1.n363 VB1.n349 0.114786
R4401 VB1.n367 VB1.n349 0.114786
R4402 VB1.n368 VB1.n348 0.114786
R4403 VB1.n372 VB1.n348 0.114786
R4404 VB1.n406 VB1.n400 0.114786
R4405 VB1.n402 VB1.n400 0.114786
R4406 VB1.n380 VB1.n378 0.114786
R4407 VB1.n384 VB1.n378 0.114786
R4408 VB1.n385 VB1.n377 0.114786
R4409 VB1.n389 VB1.n377 0.114786
R4410 VB1.n390 VB1.n376 0.114786
R4411 VB1.n394 VB1.n376 0.114786
R4412 VB1.n395 VB1.n375 0.114786
R4413 VB1.n399 VB1.n375 0.114786
R4414 VB1.n483 VB1.n477 0.114786
R4415 VB1.n479 VB1.n477 0.114786
R4416 VB1.n500 VB1.n494 0.114786
R4417 VB1.n496 VB1.n494 0.114786
R4418 VB1.n526 VB1.n489 0.114786
R4419 VB1.n522 VB1.n489 0.114786
R4420 VB1.n521 VB1.n490 0.114786
R4421 VB1.n517 VB1.n490 0.114786
R4422 VB1.n516 VB1.n491 0.114786
R4423 VB1.n512 VB1.n491 0.114786
R4424 VB1.n511 VB1.n492 0.114786
R4425 VB1.n507 VB1.n492 0.114786
R4426 VB1.n506 VB1.n493 0.114786
R4427 VB1.n502 VB1.n493 0.114786
R4428 VB1.n532 VB1.n488 0.114786
R4429 VB1.n536 VB1.n488 0.114786
R4430 VB1.n537 VB1.n487 0.114786
R4431 VB1.n541 VB1.n487 0.114786
R4432 VB1.n542 VB1.n486 0.114786
R4433 VB1.n546 VB1.n486 0.114786
R4434 VB1.n547 VB1.n485 0.114786
R4435 VB1.n551 VB1.n485 0.114786
R4436 VB1.n552 VB1.n484 0.114786
R4437 VB1.n556 VB1.n484 0.114786
R4438 VB1.n448 VB1.n442 0.114786
R4439 VB1.n444 VB1.n442 0.114786
R4440 VB1.n454 VB1.n452 0.114786
R4441 VB1.n458 VB1.n452 0.114786
R4442 VB1.n459 VB1.n451 0.114786
R4443 VB1.n463 VB1.n451 0.114786
R4444 VB1.n464 VB1.n450 0.114786
R4445 VB1.n468 VB1.n450 0.114786
R4446 VB1.n469 VB1.n449 0.114786
R4447 VB1.n473 VB1.n449 0.114786
R4448 VB1.n440 VB1.n434 0.114786
R4449 VB1.n436 VB1.n434 0.114786
R4450 VB1.n414 VB1.n412 0.114786
R4451 VB1.n418 VB1.n412 0.114786
R4452 VB1.n419 VB1.n411 0.114786
R4453 VB1.n423 VB1.n411 0.114786
R4454 VB1.n424 VB1.n410 0.114786
R4455 VB1.n428 VB1.n410 0.114786
R4456 VB1.n429 VB1.n409 0.114786
R4457 VB1.n433 VB1.n409 0.114786
R4458 VB1.n33 VB1 0.0929333
R4459 VB1.n258 VB1.n244 0.0847867
R4460 VB1.n340 VB1.n326 0.0847867
R4461 VB1 VB1.n558 0.07617
R4462 VB1.n39 VB1.n38 0.0611061
R4463 VB1.n38 VB1.n37 0.0611061
R4464 VB1.n63 VB1.n62 0.0611061
R4465 VB1.n64 VB1.n63 0.0611061
R4466 VB1.n58 VB1.n57 0.0611061
R4467 VB1.n59 VB1.n58 0.0611061
R4468 VB1.n53 VB1.n52 0.0611061
R4469 VB1.n54 VB1.n53 0.0611061
R4470 VB1.n48 VB1.n47 0.0611061
R4471 VB1.n49 VB1.n48 0.0611061
R4472 VB1.n107 VB1.n106 0.0611061
R4473 VB1.n106 VB1.n105 0.0611061
R4474 VB1.n131 VB1.n130 0.0611061
R4475 VB1.n132 VB1.n131 0.0611061
R4476 VB1.n126 VB1.n125 0.0611061
R4477 VB1.n127 VB1.n126 0.0611061
R4478 VB1.n121 VB1.n120 0.0611061
R4479 VB1.n122 VB1.n121 0.0611061
R4480 VB1.n116 VB1.n115 0.0611061
R4481 VB1.n117 VB1.n116 0.0611061
R4482 VB1.n166 VB1.n165 0.0611061
R4483 VB1.n165 VB1.n164 0.0611061
R4484 VB1.n158 VB1.n157 0.0611061
R4485 VB1.n159 VB1.n158 0.0611061
R4486 VB1.n153 VB1.n152 0.0611061
R4487 VB1.n154 VB1.n153 0.0611061
R4488 VB1.n148 VB1.n147 0.0611061
R4489 VB1.n149 VB1.n148 0.0611061
R4490 VB1.n143 VB1.n142 0.0611061
R4491 VB1.n144 VB1.n143 0.0611061
R4492 VB1.n182 VB1.n181 0.0611061
R4493 VB1.n181 VB1.n180 0.0611061
R4494 VB1.n206 VB1.n205 0.0611061
R4495 VB1.n207 VB1.n206 0.0611061
R4496 VB1.n201 VB1.n200 0.0611061
R4497 VB1.n202 VB1.n201 0.0611061
R4498 VB1.n196 VB1.n195 0.0611061
R4499 VB1.n197 VB1.n196 0.0611061
R4500 VB1.n191 VB1.n190 0.0611061
R4501 VB1.n192 VB1.n191 0.0611061
R4502 VB1.n241 VB1.n240 0.0611061
R4503 VB1.n240 VB1.n239 0.0611061
R4504 VB1.n233 VB1.n232 0.0611061
R4505 VB1.n234 VB1.n233 0.0611061
R4506 VB1.n228 VB1.n227 0.0611061
R4507 VB1.n229 VB1.n228 0.0611061
R4508 VB1.n223 VB1.n222 0.0611061
R4509 VB1.n224 VB1.n223 0.0611061
R4510 VB1.n218 VB1.n217 0.0611061
R4511 VB1.n219 VB1.n218 0.0611061
R4512 VB1.n323 VB1.n322 0.0611061
R4513 VB1.n322 VB1.n321 0.0611061
R4514 VB1.n315 VB1.n314 0.0611061
R4515 VB1.n316 VB1.n315 0.0611061
R4516 VB1.n310 VB1.n309 0.0611061
R4517 VB1.n311 VB1.n310 0.0611061
R4518 VB1.n305 VB1.n304 0.0611061
R4519 VB1.n306 VB1.n305 0.0611061
R4520 VB1.n300 VB1.n299 0.0611061
R4521 VB1.n301 VB1.n300 0.0611061
R4522 VB1.n346 VB1.n345 0.0611061
R4523 VB1.n345 VB1.n344 0.0611061
R4524 VB1.n370 VB1.n369 0.0611061
R4525 VB1.n371 VB1.n370 0.0611061
R4526 VB1.n365 VB1.n364 0.0611061
R4527 VB1.n366 VB1.n365 0.0611061
R4528 VB1.n360 VB1.n359 0.0611061
R4529 VB1.n361 VB1.n360 0.0611061
R4530 VB1.n355 VB1.n354 0.0611061
R4531 VB1.n356 VB1.n355 0.0611061
R4532 VB1.n482 VB1.n481 0.0611061
R4533 VB1.n481 VB1.n480 0.0611061
R4534 VB1.n554 VB1.n553 0.0611061
R4535 VB1.n555 VB1.n554 0.0611061
R4536 VB1.n549 VB1.n548 0.0611061
R4537 VB1.n550 VB1.n549 0.0611061
R4538 VB1.n544 VB1.n543 0.0611061
R4539 VB1.n545 VB1.n544 0.0611061
R4540 VB1.n539 VB1.n538 0.0611061
R4541 VB1.n540 VB1.n539 0.0611061
R4542 VB1.n534 VB1.n533 0.0611061
R4543 VB1.n535 VB1.n534 0.0611061
R4544 VB1.n447 VB1.n446 0.0611061
R4545 VB1.n446 VB1.n445 0.0611061
R4546 VB1.n471 VB1.n470 0.0611061
R4547 VB1.n472 VB1.n471 0.0611061
R4548 VB1.n466 VB1.n465 0.0611061
R4549 VB1.n467 VB1.n466 0.0611061
R4550 VB1.n461 VB1.n460 0.0611061
R4551 VB1.n462 VB1.n461 0.0611061
R4552 VB1.n456 VB1.n455 0.0611061
R4553 VB1.n457 VB1.n456 0.0611061
R4554 VB1.n30 VB1.n29 0.0605379
R4555 VB1.n22 VB1.n21 0.0605379
R4556 VB1.n17 VB1.n16 0.0605379
R4557 VB1.n12 VB1.n11 0.0605379
R4558 VB1.n7 VB1.n6 0.0605379
R4559 VB1.n98 VB1.n97 0.0605379
R4560 VB1.n90 VB1.n89 0.0605379
R4561 VB1.n85 VB1.n84 0.0605379
R4562 VB1.n80 VB1.n79 0.0605379
R4563 VB1.n75 VB1.n74 0.0605379
R4564 VB1.n405 VB1.n404 0.0605379
R4565 VB1.n397 VB1.n396 0.0605379
R4566 VB1.n392 VB1.n391 0.0605379
R4567 VB1.n387 VB1.n386 0.0605379
R4568 VB1.n382 VB1.n381 0.0605379
R4569 VB1.n505 VB1.n504 0.0605379
R4570 VB1.n510 VB1.n509 0.0605379
R4571 VB1.n515 VB1.n514 0.0605379
R4572 VB1.n520 VB1.n519 0.0605379
R4573 VB1.n525 VB1.n524 0.0605379
R4574 VB1.n499 VB1.n498 0.0605379
R4575 VB1.n439 VB1.n438 0.0605379
R4576 VB1.n431 VB1.n430 0.0605379
R4577 VB1.n426 VB1.n425 0.0605379
R4578 VB1.n421 VB1.n420 0.0605379
R4579 VB1.n416 VB1.n415 0.0605379
R4580 VB1.n29 VB1.n28 0.0603695
R4581 VB1.n23 VB1.n22 0.0603695
R4582 VB1.n18 VB1.n17 0.0603695
R4583 VB1.n13 VB1.n12 0.0603695
R4584 VB1.n8 VB1.n7 0.0603695
R4585 VB1.n97 VB1.n96 0.0603695
R4586 VB1.n91 VB1.n90 0.0603695
R4587 VB1.n86 VB1.n85 0.0603695
R4588 VB1.n81 VB1.n80 0.0603695
R4589 VB1.n76 VB1.n75 0.0603695
R4590 VB1.n404 VB1.n403 0.0603695
R4591 VB1.n398 VB1.n397 0.0603695
R4592 VB1.n393 VB1.n392 0.0603695
R4593 VB1.n388 VB1.n387 0.0603695
R4594 VB1.n383 VB1.n382 0.0603695
R4595 VB1.n504 VB1.n503 0.0603695
R4596 VB1.n509 VB1.n508 0.0603695
R4597 VB1.n514 VB1.n513 0.0603695
R4598 VB1.n519 VB1.n518 0.0603695
R4599 VB1.n524 VB1.n523 0.0603695
R4600 VB1.n498 VB1.n497 0.0603695
R4601 VB1.n438 VB1.n437 0.0603695
R4602 VB1.n432 VB1.n431 0.0603695
R4603 VB1.n427 VB1.n426 0.0603695
R4604 VB1.n422 VB1.n421 0.0603695
R4605 VB1.n417 VB1.n416 0.0603695
R4606 VB1.n264 VB1.n263 0.0603541
R4607 VB1.n288 VB1.n287 0.0603541
R4608 VB1.n283 VB1.n282 0.0603541
R4609 VB1.n278 VB1.n277 0.0603541
R4610 VB1.n273 VB1.n272 0.0603541
R4611 VB1.n263 VB1.n262 0.0601312
R4612 VB1.n289 VB1.n288 0.0601312
R4613 VB1.n284 VB1.n283 0.0601312
R4614 VB1.n279 VB1.n278 0.0601312
R4615 VB1.n274 VB1.n273 0.0601312
R4616 VB1.n292 VB1.n258 0.0594067
R4617 VB1.n374 VB1.n340 0.0589367
R4618 VB1.n210 VB1.n176 0.05831
R4619 VB1.n326 VB1.n292 0.0288567
R4620 VB1.n169 VB1.n135 0.0287
R4621 VB1.n244 VB1.n210 0.0287
R4622 VB1.n101 VB1.n67 0.0271333
R4623 VB1.n408 VB1.n374 0.0271333
R4624 VB1.n558 VB1.n476 0.0271333
R4625 AVDD.n295 AVDD.n294 20442.4
R4626 AVDD.n1734 AVDD.n1733 20442.4
R4627 AVDD.n2997 AVDD.n298 2180.52
R4628 AVDD.n3109 AVDD.n3108 2180.52
R4629 AVDD.n1137 AVDD.n200 1160.36
R4630 AVDD.n498 AVDD.n497 1150.59
R4631 AVDD.n1892 AVDD.n503 1083.53
R4632 AVDD.n2185 AVDD.n92 1002.35
R4633 AVDD.n978 AVDD.n775 949.413
R4634 AVDD.n3295 AVDD.n97 935.294
R4635 AVDD.n976 AVDD.n778 896.471
R4636 AVDD.n3122 AVDD.n3121 850.588
R4637 AVDD.n1138 AVDD.n593 847.059
R4638 AVDD.n1135 AVDD.n682 794.119
R4639 AVDD.n2992 AVDD.n2991 240
R4640 AVDD.n2989 AVDD.n306 240
R4641 AVDD.n2979 AVDD.n318 240
R4642 AVDD.n2977 AVDD.n319 240
R4643 AVDD.n2970 AVDD.n2969 240
R4644 AVDD.n2967 AVDD.n325 240
R4645 AVDD.n2960 AVDD.n2959 240
R4646 AVDD.n2957 AVDD.n334 240
R4647 AVDD.n2950 AVDD.n2949 240
R4648 AVDD.n2947 AVDD.n342 240
R4649 AVDD.n2940 AVDD.n357 240
R4650 AVDD.n2938 AVDD.n358 240
R4651 AVDD.n2930 AVDD.n2929 240
R4652 AVDD.n2927 AVDD.n364 240
R4653 AVDD.n2920 AVDD.n2919 240
R4654 AVDD.n2917 AVDD.n378 240
R4655 AVDD.n2910 AVDD.n2909 240
R4656 AVDD.n2907 AVDD.n400 240
R4657 AVDD.n2900 AVDD.n2899 240
R4658 AVDD.n2897 AVDD.n409 240
R4659 AVDD.n2886 AVDD.n2885 240
R4660 AVDD.n2883 AVDD.n417 240
R4661 AVDD.n2876 AVDD.n2875 240
R4662 AVDD.n2873 AVDD.n426 240
R4663 AVDD.n2863 AVDD.n440 240
R4664 AVDD.n2861 AVDD.n441 240
R4665 AVDD.n2854 AVDD.n2853 240
R4666 AVDD.n2851 AVDD.n447 240
R4667 AVDD.n2844 AVDD.n455 240
R4668 AVDD.n2842 AVDD.n456 240
R4669 AVDD.n1923 AVDD.n498 240
R4670 AVDD.n1923 AVDD.n500 240
R4671 AVDD.n1903 AVDD.n500 240
R4672 AVDD.n1903 AVDD.n1900 240
R4673 AVDD.n1911 AVDD.n1900 240
R4674 AVDD.n1913 AVDD.n1911 240
R4675 AVDD.n1913 AVDD.n481 240
R4676 AVDD.n1930 AVDD.n481 240
R4677 AVDD.n1930 AVDD.n469 240
R4678 AVDD.n2831 AVDD.n469 240
R4679 AVDD.n2831 AVDD.n470 240
R4680 AVDD.n1942 AVDD.n470 240
R4681 AVDD.n1943 AVDD.n1942 240
R4682 AVDD.n1944 AVDD.n1943 240
R4683 AVDD.n2408 AVDD.n1944 240
R4684 AVDD.n2408 AVDD.n2407 240
R4685 AVDD.n2407 AVDD.n2402 240
R4686 AVDD.n2402 AVDD.n1962 240
R4687 AVDD.n1963 AVDD.n1962 240
R4688 AVDD.n1964 AVDD.n1963 240
R4689 AVDD.n2375 AVDD.n1964 240
R4690 AVDD.n2375 AVDD.n1979 240
R4691 AVDD.n1980 AVDD.n1979 240
R4692 AVDD.n1982 AVDD.n1980 240
R4693 AVDD.n2440 AVDD.n1982 240
R4694 AVDD.n2440 AVDD.n1993 240
R4695 AVDD.n1994 AVDD.n1993 240
R4696 AVDD.n1995 AVDD.n1994 240
R4697 AVDD.n2517 AVDD.n1995 240
R4698 AVDD.n2517 AVDD.n2006 240
R4699 AVDD.n2007 AVDD.n2006 240
R4700 AVDD.n2008 AVDD.n2007 240
R4701 AVDD.n2462 AVDD.n2008 240
R4702 AVDD.n2468 AVDD.n2462 240
R4703 AVDD.n2469 AVDD.n2468 240
R4704 AVDD.n2469 AVDD.n2026 240
R4705 AVDD.n2027 AVDD.n2026 240
R4706 AVDD.n2028 AVDD.n2027 240
R4707 AVDD.n2479 AVDD.n2028 240
R4708 AVDD.n2479 AVDD.n2038 240
R4709 AVDD.n2039 AVDD.n2038 240
R4710 AVDD.n2040 AVDD.n2039 240
R4711 AVDD.n2365 AVDD.n2040 240
R4712 AVDD.n2365 AVDD.n2052 240
R4713 AVDD.n2053 AVDD.n2052 240
R4714 AVDD.n2054 AVDD.n2053 240
R4715 AVDD.n2542 AVDD.n2054 240
R4716 AVDD.n2542 AVDD.n2075 240
R4717 AVDD.n2076 AVDD.n2075 240
R4718 AVDD.n2077 AVDD.n2076 240
R4719 AVDD.n2556 AVDD.n2077 240
R4720 AVDD.n2557 AVDD.n2556 240
R4721 AVDD.n2557 AVDD.n2093 240
R4722 AVDD.n2094 AVDD.n2093 240
R4723 AVDD.n2095 AVDD.n2094 240
R4724 AVDD.n2568 AVDD.n2095 240
R4725 AVDD.n2568 AVDD.n2567 240
R4726 AVDD.n2567 AVDD.n2111 240
R4727 AVDD.n2112 AVDD.n2111 240
R4728 AVDD.n2113 AVDD.n2112 240
R4729 AVDD.n2593 AVDD.n2113 240
R4730 AVDD.n2593 AVDD.n2125 240
R4731 AVDD.n2126 AVDD.n2125 240
R4732 AVDD.n2127 AVDD.n2126 240
R4733 AVDD.n2608 AVDD.n2127 240
R4734 AVDD.n2608 AVDD.n2144 240
R4735 AVDD.n2145 AVDD.n2144 240
R4736 AVDD.n2146 AVDD.n2145 240
R4737 AVDD.n2622 AVDD.n2146 240
R4738 AVDD.n2623 AVDD.n2622 240
R4739 AVDD.n2623 AVDD.n2162 240
R4740 AVDD.n2163 AVDD.n2162 240
R4741 AVDD.n2164 AVDD.n2163 240
R4742 AVDD.n2197 AVDD.n2164 240
R4743 AVDD.n2208 AVDD.n2197 240
R4744 AVDD.n2208 AVDD.n2201 240
R4745 AVDD.n2201 AVDD.n2199 240
R4746 AVDD.n2199 AVDD.n2183 240
R4747 AVDD.n2184 AVDD.n2183 240
R4748 AVDD.n2640 AVDD.n2184 240
R4749 AVDD.n2640 AVDD.n2185 240
R4750 AVDD.n1333 AVDD.n94 240
R4751 AVDD.n1348 AVDD.n1347 240
R4752 AVDD.n1352 AVDD.n1351 240
R4753 AVDD.n1361 AVDD.n1360 240
R4754 AVDD.n1365 AVDD.n1364 240
R4755 AVDD.n1374 AVDD.n1373 240
R4756 AVDD.n1378 AVDD.n1377 240
R4757 AVDD.n1389 AVDD.n1388 240
R4758 AVDD.n1698 AVDD.n1697 240
R4759 AVDD.n1690 AVDD.n1689 240
R4760 AVDD.n1679 AVDD.n1678 240
R4761 AVDD.n1672 AVDD.n1671 240
R4762 AVDD.n1668 AVDD.n1667 240
R4763 AVDD.n1659 AVDD.n1658 240
R4764 AVDD.n1655 AVDD.n1654 240
R4765 AVDD.n1647 AVDD.n1646 240
R4766 AVDD.n1640 AVDD.n1639 240
R4767 AVDD.n1636 AVDD.n1635 240
R4768 AVDD.n1624 AVDD.n1623 240
R4769 AVDD.n1443 AVDD.n62 240
R4770 AVDD.n1613 AVDD.n93 240
R4771 AVDD.n1450 AVDD.n1449 240
R4772 AVDD.n1607 AVDD.n1606 240
R4773 AVDD.n1599 AVDD.n1598 240
R4774 AVDD.n1595 AVDD.n1594 240
R4775 AVDD.n1587 AVDD.n1586 240
R4776 AVDD.n1580 AVDD.n1579 240
R4777 AVDD.n1576 AVDD.n1575 240
R4778 AVDD.n1568 AVDD.n1567 240
R4779 AVDD.n1557 AVDD.n1556 240
R4780 AVDD.n1501 AVDD.n1500 240
R4781 AVDD.n1550 AVDD.n1549 240
R4782 AVDD.n1541 AVDD.n1540 240
R4783 AVDD.n1537 AVDD.n1536 240
R4784 AVDD.n1529 AVDD.n1528 240
R4785 AVDD.n1525 AVDD.n1524 240
R4786 AVDD.n1518 AVDD.n12 240
R4787 AVDD.n3299 AVDD.n11 240
R4788 AVDD.n2240 AVDD.n2239 240
R4789 AVDD.n2243 AVDD.n2242 240
R4790 AVDD.n2255 AVDD.n2254 240
R4791 AVDD.n2265 AVDD.n2264 240
R4792 AVDD.n2269 AVDD.n2268 240
R4793 AVDD.n2276 AVDD.n2275 240
R4794 AVDD.n2291 AVDD.n2290 240
R4795 AVDD.n2295 AVDD.n2294 240
R4796 AVDD.n2304 AVDD.n2303 240
R4797 AVDD.n2308 AVDD.n2307 240
R4798 AVDD.n2316 AVDD.n2315 240
R4799 AVDD.n2328 AVDD.n2327 240
R4800 AVDD.n2324 AVDD.n92 240
R4801 AVDD.n1921 AVDD.n503 240
R4802 AVDD.n1921 AVDD.n504 240
R4803 AVDD.n1906 AVDD.n504 240
R4804 AVDD.n1908 AVDD.n1906 240
R4805 AVDD.n1908 AVDD.n1898 240
R4806 AVDD.n1915 AVDD.n1898 240
R4807 AVDD.n1915 AVDD.n479 240
R4808 AVDD.n1932 AVDD.n479 240
R4809 AVDD.n1932 AVDD.n473 240
R4810 AVDD.n2829 AVDD.n473 240
R4811 AVDD.n2829 AVDD.n474 240
R4812 AVDD.n2822 AVDD.n474 240
R4813 AVDD.n2822 AVDD.n1941 240
R4814 AVDD.n2818 AVDD.n1941 240
R4815 AVDD.n2818 AVDD.n1946 240
R4816 AVDD.n2405 AVDD.n1946 240
R4817 AVDD.n2405 AVDD.n1959 240
R4818 AVDD.n2808 AVDD.n1959 240
R4819 AVDD.n2808 AVDD.n1960 240
R4820 AVDD.n2804 AVDD.n1960 240
R4821 AVDD.n2804 AVDD.n1965 240
R4822 AVDD.n2795 AVDD.n1965 240
R4823 AVDD.n2795 AVDD.n1977 240
R4824 AVDD.n2792 AVDD.n1977 240
R4825 AVDD.n2792 AVDD.n1983 240
R4826 AVDD.n2783 AVDD.n1983 240
R4827 AVDD.n2783 AVDD.n1992 240
R4828 AVDD.n2779 AVDD.n1992 240
R4829 AVDD.n2779 AVDD.n1997 240
R4830 AVDD.n2771 AVDD.n1997 240
R4831 AVDD.n2771 AVDD.n2005 240
R4832 AVDD.n2767 AVDD.n2005 240
R4833 AVDD.n2767 AVDD.n2010 240
R4834 AVDD.n2466 AVDD.n2010 240
R4835 AVDD.n2466 AVDD.n2023 240
R4836 AVDD.n2757 AVDD.n2023 240
R4837 AVDD.n2757 AVDD.n2024 240
R4838 AVDD.n2753 AVDD.n2024 240
R4839 AVDD.n2753 AVDD.n2029 240
R4840 AVDD.n2744 AVDD.n2029 240
R4841 AVDD.n2744 AVDD.n2036 240
R4842 AVDD.n2740 AVDD.n2036 240
R4843 AVDD.n2740 AVDD.n2041 240
R4844 AVDD.n2731 AVDD.n2041 240
R4845 AVDD.n2731 AVDD.n2050 240
R4846 AVDD.n2727 AVDD.n2050 240
R4847 AVDD.n2727 AVDD.n2056 240
R4848 AVDD.n2719 AVDD.n2056 240
R4849 AVDD.n2719 AVDD.n2074 240
R4850 AVDD.n2715 AVDD.n2074 240
R4851 AVDD.n2715 AVDD.n2079 240
R4852 AVDD.n2090 AVDD.n2079 240
R4853 AVDD.n2707 AVDD.n2090 240
R4854 AVDD.n2707 AVDD.n2091 240
R4855 AVDD.n2703 AVDD.n2091 240
R4856 AVDD.n2703 AVDD.n2097 240
R4857 AVDD.n2108 AVDD.n2097 240
R4858 AVDD.n2693 AVDD.n2108 240
R4859 AVDD.n2693 AVDD.n2109 240
R4860 AVDD.n2689 AVDD.n2109 240
R4861 AVDD.n2689 AVDD.n2114 240
R4862 AVDD.n2680 AVDD.n2114 240
R4863 AVDD.n2680 AVDD.n2123 240
R4864 AVDD.n2676 AVDD.n2123 240
R4865 AVDD.n2676 AVDD.n2129 240
R4866 AVDD.n2668 AVDD.n2129 240
R4867 AVDD.n2668 AVDD.n2143 240
R4868 AVDD.n2664 AVDD.n2143 240
R4869 AVDD.n2664 AVDD.n2148 240
R4870 AVDD.n2159 AVDD.n2148 240
R4871 AVDD.n2656 AVDD.n2159 240
R4872 AVDD.n2656 AVDD.n2160 240
R4873 AVDD.n2652 AVDD.n2160 240
R4874 AVDD.n2652 AVDD.n2166 240
R4875 AVDD.n2206 AVDD.n2166 240
R4876 AVDD.n2206 AVDD.n2204 240
R4877 AVDD.n2204 AVDD.n2179 240
R4878 AVDD.n2646 AVDD.n2179 240
R4879 AVDD.n2646 AVDD.n2181 240
R4880 AVDD.n2642 AVDD.n2181 240
R4881 AVDD.n2642 AVDD.n97 240
R4882 AVDD.n1890 AVDD.n513 240
R4883 AVDD.n1879 AVDD.n1878 240
R4884 AVDD.n1876 AVDD.n522 240
R4885 AVDD.n1869 AVDD.n531 240
R4886 AVDD.n1867 AVDD.n532 240
R4887 AVDD.n1857 AVDD.n544 240
R4888 AVDD.n1855 AVDD.n545 240
R4889 AVDD.n1848 AVDD.n1847 240
R4890 AVDD.n1845 AVDD.n551 240
R4891 AVDD.n1837 AVDD.n1836 240
R4892 AVDD.n1834 AVDD.n1146 240
R4893 AVDD.n1824 AVDD.n1159 240
R4894 AVDD.n1822 AVDD.n1821 240
R4895 AVDD.n1819 AVDD.n1162 240
R4896 AVDD.n1812 AVDD.n1811 240
R4897 AVDD.n1809 AVDD.n1171 240
R4898 AVDD.n1799 AVDD.n1185 240
R4899 AVDD.n1797 AVDD.n1186 240
R4900 AVDD.n1790 AVDD.n1789 240
R4901 AVDD.n1787 AVDD.n1192 240
R4902 AVDD.n1780 AVDD.n1779 240
R4903 AVDD.n1777 AVDD.n1201 240
R4904 AVDD.n1770 AVDD.n1769 240
R4905 AVDD.n1767 AVDD.n1207 240
R4906 AVDD.n1759 AVDD.n1758 240
R4907 AVDD.n1756 AVDD.n1221 240
R4908 AVDD.n1748 AVDD.n1747 240
R4909 AVDD.n1745 AVDD.n1229 240
R4910 AVDD.n1738 AVDD.n1737 240
R4911 AVDD.n3103 AVDD.n3102 240
R4912 AVDD.n3100 AVDD.n201 240
R4913 AVDD.n3093 AVDD.n3092 240
R4914 AVDD.n3090 AVDD.n215 240
R4915 AVDD.n3083 AVDD.n3082 240
R4916 AVDD.n3080 AVDD.n222 240
R4917 AVDD.n3070 AVDD.n236 240
R4918 AVDD.n3068 AVDD.n237 240
R4919 AVDD.n3061 AVDD.n3060 240
R4920 AVDD.n3058 AVDD.n244 240
R4921 AVDD.n3047 AVDD.n3046 240
R4922 AVDD.n3044 AVDD.n254 240
R4923 AVDD.n3037 AVDD.n263 240
R4924 AVDD.n3035 AVDD.n264 240
R4925 AVDD.n3025 AVDD.n276 240
R4926 AVDD.n3023 AVDD.n277 240
R4927 AVDD.n3016 AVDD.n3015 240
R4928 AVDD.n3013 AVDD.n284 240
R4929 AVDD.n3002 AVDD.n3001 240
R4930 AVDD.n96 AVDD.n95 240
R4931 AVDD.n3285 AVDD.n95 240
R4932 AVDD.n3279 AVDD.n3278 240
R4933 AVDD.n3275 AVDD.n3274 240
R4934 AVDD.n3266 AVDD.n3265 240
R4935 AVDD.n3262 AVDD.n3261 240
R4936 AVDD.n3254 AVDD.n3253 240
R4937 AVDD.n3250 AVDD.n3249 240
R4938 AVDD.n3242 AVDD.n3241 240
R4939 AVDD.n3235 AVDD.n3234 240
R4940 AVDD.n3231 AVDD.n3230 240
R4941 AVDD.n138 AVDD.n137 240
R4942 AVDD.n3220 AVDD.n3219 240
R4943 AVDD.n3215 AVDD.n3214 240
R4944 AVDD.n3207 AVDD.n3206 240
R4945 AVDD.n3203 AVDD.n3202 240
R4946 AVDD.n156 AVDD.n155 240
R4947 AVDD.n3192 AVDD.n3191 240
R4948 AVDD.n3184 AVDD.n3183 240
R4949 AVDD.n3180 AVDD.n3179 240
R4950 AVDD.n3172 AVDD.n3171 240
R4951 AVDD.n3168 AVDD.n3167 240
R4952 AVDD.n3160 AVDD.n3159 240
R4953 AVDD.n3149 AVDD.n3148 240
R4954 AVDD.n3145 AVDD.n3144 240
R4955 AVDD.n3137 AVDD.n3136 240
R4956 AVDD.n3133 AVDD.n3132 240
R4957 AVDD.n3118 AVDD.n3117 240
R4958 AVDD.n187 AVDD.n42 240
R4959 AVDD.n976 AVDD.n769 240
R4960 AVDD.n987 AVDD.n769 240
R4961 AVDD.n987 AVDD.n764 240
R4962 AVDD.n998 AVDD.n764 240
R4963 AVDD.n998 AVDD.n755 240
R4964 AVDD.n1022 AVDD.n755 240
R4965 AVDD.n1022 AVDD.n751 240
R4966 AVDD.n1033 AVDD.n751 240
R4967 AVDD.n1033 AVDD.n739 240
R4968 AVDD.n1063 AVDD.n739 240
R4969 AVDD.n1063 AVDD.n740 240
R4970 AVDD.n1059 AVDD.n740 240
R4971 AVDD.n1059 AVDD.n731 240
R4972 AVDD.n1077 AVDD.n731 240
R4973 AVDD.n1077 AVDD.n719 240
R4974 AVDD.n1095 AVDD.n719 240
R4975 AVDD.n1095 AVDD.n720 240
R4976 AVDD.n720 AVDD.n706 240
R4977 AVDD.n1112 AVDD.n706 240
R4978 AVDD.n1113 AVDD.n1112 240
R4979 AVDD.n1113 AVDD.n687 240
R4980 AVDD.n1124 AVDD.n687 240
R4981 AVDD.n1125 AVDD.n1124 240
R4982 AVDD.n1125 AVDD.n682 240
R4983 AVDD.n681 AVDD.n679 240
R4984 AVDD.n679 AVDD.n677 240
R4985 AVDD.n599 AVDD.n597 240
R4986 AVDD.n604 AVDD.n602 240
R4987 AVDD.n609 AVDD.n607 240
R4988 AVDD.n614 AVDD.n613 240
R4989 AVDD.n619 AVDD.n617 240
R4990 AVDD.n624 AVDD.n622 240
R4991 AVDD.n629 AVDD.n627 240
R4992 AVDD.n634 AVDD.n632 240
R4993 AVDD.n639 AVDD.n637 240
R4994 AVDD.n644 AVDD.n642 240
R4995 AVDD.n649 AVDD.n647 240
R4996 AVDD.n654 AVDD.n652 240
R4997 AVDD.n659 AVDD.n658 240
R4998 AVDD.n664 AVDD.n662 240
R4999 AVDD.n669 AVDD.n667 240
R5000 AVDD.n674 AVDD.n672 240
R5001 AVDD.n1138 AVDD.n592 240
R5002 AVDD.n978 AVDD.n770 240
R5003 AVDD.n985 AVDD.n770 240
R5004 AVDD.n985 AVDD.n762 240
R5005 AVDD.n1000 AVDD.n762 240
R5006 AVDD.n1000 AVDD.n757 240
R5007 AVDD.n1019 AVDD.n757 240
R5008 AVDD.n1019 AVDD.n749 240
R5009 AVDD.n1035 AVDD.n749 240
R5010 AVDD.n1036 AVDD.n1035 240
R5011 AVDD.n1036 AVDD.n742 240
R5012 AVDD.n743 AVDD.n742 240
R5013 AVDD.n1050 AVDD.n743 240
R5014 AVDD.n1050 AVDD.n744 240
R5015 AVDD.n744 AVDD.n729 240
R5016 AVDD.n1080 AVDD.n729 240
R5017 AVDD.n1080 AVDD.n721 240
R5018 AVDD.n1092 AVDD.n721 240
R5019 AVDD.n1092 AVDD.n709 240
R5020 AVDD.n1110 AVDD.n709 240
R5021 AVDD.n1110 AVDD.n690 240
R5022 AVDD.n1121 AVDD.n690 240
R5023 AVDD.n1121 AVDD.n686 240
R5024 AVDD.n1127 AVDD.n686 240
R5025 AVDD.n1127 AVDD.n593 240
R5026 AVDD.n960 AVDD.n952 240
R5027 AVDD.n963 AVDD.n962 240
R5028 AVDD.n965 AVDD.n949 240
R5029 AVDD.n940 AVDD.n791 240
R5030 AVDD.n938 AVDD.n792 240
R5031 AVDD.n931 AVDD.n929 240
R5032 AVDD.n927 AVDD.n797 240
R5033 AVDD.n918 AVDD.n916 240
R5034 AVDD.n909 AVDD.n809 240
R5035 AVDD.n907 AVDD.n810 240
R5036 AVDD.n899 AVDD.n897 240
R5037 AVDD.n890 AVDD.n823 240
R5038 AVDD.n888 AVDD.n824 240
R5039 AVDD.n881 AVDD.n879 240
R5040 AVDD.n868 AVDD.n867 240
R5041 AVDD.n870 AVDD.n866 240
R5042 AVDD.n859 AVDD.n844 240
R5043 AVDD.n857 AVDD.n846 240
R5044 AVDD.n1252 AVDD.t24 232.707
R5045 AVDD.n1249 AVDD.t124 232.707
R5046 AVDD.n1251 AVDD.t61 232.707
R5047 AVDD.n1257 AVDD.t88 232.707
R5048 AVDD.n1266 AVDD.t76 232.707
R5049 AVDD.n1277 AVDD.t106 232.707
R5050 AVDD.n1274 AVDD.t93 232.707
R5051 AVDD.n1276 AVDD.t28 232.707
R5052 AVDD.n1282 AVDD.t12 232.707
R5053 AVDD.n1291 AVDD.t47 232.707
R5054 AVDD.n1468 AVDD.t73 232.707
R5055 AVDD.n1465 AVDD.t57 232.707
R5056 AVDD.n1467 AVDD.t92 232.707
R5057 AVDD.n1473 AVDD.t13 232.707
R5058 AVDD.n1482 AVDD.t109 232.707
R5059 AVDD.n382 AVDD.t77 232.707
R5060 AVDD.n3 AVDD.t9 232.707
R5061 AVDD.n384 AVDD.t40 232.707
R5062 AVDD.n385 AVDD.t116 232.707
R5063 AVDD.n6 AVDD.t70 232.707
R5064 AVDD.n2337 AVDD.t112 232.703
R5065 AVDD.n2578 AVDD.t68 232.703
R5066 AVDD.n2370 AVDD.t60 232.703
R5067 AVDD.n2444 AVDD.t83 232.703
R5068 AVDD.n2387 AVDD.t121 232.703
R5069 AVDD.n1252 AVDD.t78 232.703
R5070 AVDD.n1249 AVDD.t65 232.703
R5071 AVDD.n1251 AVDD.t102 232.703
R5072 AVDD.n1257 AVDD.t31 232.703
R5073 AVDD.n1266 AVDD.t118 232.703
R5074 AVDD.n1277 AVDD.t59 232.703
R5075 AVDD.n1274 AVDD.t44 232.703
R5076 AVDD.n1276 AVDD.t82 232.703
R5077 AVDD.n1282 AVDD.t126 232.703
R5078 AVDD.n1291 AVDD.t96 232.703
R5079 AVDD.n1724 AVDD.t100 232.703
R5080 AVDD.n1716 AVDD.t84 232.703
R5081 AVDD.n1242 AVDD.t17 232.703
R5082 AVDD.n1243 AVDD.t67 232.703
R5083 AVDD.n1709 AVDD.t39 232.703
R5084 AVDD.n1468 AVDD.t66 232.703
R5085 AVDD.n1465 AVDD.t26 232.703
R5086 AVDD.n1467 AVDD.t46 232.703
R5087 AVDD.n1473 AVDD.t108 232.703
R5088 AVDD.n1482 AVDD.t117 232.703
R5089 AVDD.n382 AVDD.t99 232.703
R5090 AVDD.n3 AVDD.t10 232.703
R5091 AVDD.n384 AVDD.t72 232.703
R5092 AVDD.n385 AVDD.t37 232.703
R5093 AVDD.n6 AVDD.t89 232.703
R5094 AVDD.n1724 AVDD.t69 232.328
R5095 AVDD.n1716 AVDD.t55 232.328
R5096 AVDD.n1242 AVDD.t90 232.328
R5097 AVDD.n1243 AVDD.t25 232.328
R5098 AVDD.n1709 AVDD.t107 232.328
R5099 AVDD.n1428 AVDD.t103 232.328
R5100 AVDD.n1411 AVDD.t14 232.327
R5101 AVDD.n1413 AVDD.t30 232.327
R5102 AVDD.n1419 AVDD.t98 232.327
R5103 AVDD.n1414 AVDD.t50 232.327
R5104 AVDD.n1300 AVDD.t119 232.317
R5105 AVDD.n1303 AVDD.t21 232.317
R5106 AVDD.n1302 AVDD.t52 232.317
R5107 AVDD.n1308 AVDD.t87 232.317
R5108 AVDD.n1317 AVDD.t75 232.317
R5109 AVDD.n713 AVDD.t6 232.169
R5110 AVDD.n714 AVDD.t7 231.998
R5111 AVDD.n1300 AVDD.t41 231.946
R5112 AVDD.n1303 AVDD.t51 231.946
R5113 AVDD.n1302 AVDD.t81 231.946
R5114 AVDD.n1308 AVDD.t125 231.946
R5115 AVDD.n1317 AVDD.t95 231.946
R5116 AVDD.n1411 AVDD.t104 231.942
R5117 AVDD.n1413 AVDD.t43 231.942
R5118 AVDD.n1419 AVDD.t79 231.942
R5119 AVDD.n1414 AVDD.t122 231.942
R5120 AVDD.n1428 AVDD.t62 231.94
R5121 AVDD.n1106 AVDD.t4 231.673
R5122 AVDD.n713 AVDD.t3 231.673
R5123 AVDD.n714 AVDD.t5 231.673
R5124 AVDD.n2337 AVDD.t390 231.644
R5125 AVDD.t254 AVDD.n2578 231.644
R5126 AVDD.n2356 AVDD.t190 231.644
R5127 AVDD.t217 AVDD.n2370 231.644
R5128 AVDD.n2444 AVDD.t295 231.644
R5129 AVDD.n2387 AVDD.t411 231.644
R5130 AVDD.n1130 AVDD.t305 231.644
R5131 AVDD.n1105 AVDD.t304 231.644
R5132 AVDD.n715 AVDD.t328 231.644
R5133 AVDD.n753 AVDD.t273 231.644
R5134 AVDD.n992 AVDD.t154 231.644
R5135 AVDD.n781 AVDD.t153 231.644
R5136 AVDD.n1088 AVDD.t259 231.644
R5137 AVDD.t173 AVDD.n1006 231.644
R5138 AVDD.n2660 AVDD.t239 231.644
R5139 AVDD.t383 AVDD.n2102 231.644
R5140 AVDD.n2711 AVDD.t139 231.644
R5141 AVDD.n2775 AVDD.t297 231.644
R5142 AVDD.n1990 AVDD.t179 231.644
R5143 AVDD.t420 AVDD.n1938 231.644
R5144 AVDD.n1130 AVDD.t351 231.643
R5145 AVDD.n1105 AVDD.t350 231.643
R5146 AVDD.n1130 AVDD.t151 231.643
R5147 AVDD.n1105 AVDD.t150 231.643
R5148 AVDD.n1130 AVDD.t184 231.643
R5149 AVDD.n1105 AVDD.t183 231.643
R5150 AVDD.n1130 AVDD.t280 231.643
R5151 AVDD.n1105 AVDD.t279 231.643
R5152 AVDD.n1130 AVDD.t414 231.643
R5153 AVDD.n1105 AVDD.t413 231.643
R5154 AVDD.n1130 AVDD.t225 231.643
R5155 AVDD.n1105 AVDD.t224 231.643
R5156 AVDD.n1885 AVDD.t325 220.367
R5157 AVDD.n1884 AVDD.t335 220.367
R5158 AVDD.n1862 AVDD.t187 220.367
R5159 AVDD.n538 AVDD.t200 220.367
R5160 AVDD.n1829 AVDD.t362 220.367
R5161 AVDD.n1153 AVDD.t379 220.367
R5162 AVDD.n1804 AVDD.t136 220.367
R5163 AVDD.n1179 AVDD.t147 220.367
R5164 AVDD.n1214 AVDD.t308 220.367
R5165 AVDD.n1213 AVDD.t310 220.367
R5166 AVDD.n1238 AVDD.t157 220.367
R5167 AVDD.n1236 AVDD.t165 220.367
R5168 AVDD.n209 AVDD.t176 220.367
R5169 AVDD.n207 AVDD.t181 220.367
R5170 AVDD.n3075 AVDD.t338 220.367
R5171 AVDD.n230 AVDD.t343 220.367
R5172 AVDD.n3053 AVDD.t160 220.367
R5173 AVDD.n3052 AVDD.t169 220.367
R5174 AVDD.n3030 AVDD.t322 220.367
R5175 AVDD.n270 AVDD.t330 220.367
R5176 AVDD.n3008 AVDD.t215 220.367
R5177 AVDD.n3007 AVDD.t284 220.367
R5178 AVDD.n2984 AVDD.t333 220.367
R5179 AVDD.n312 AVDD.t418 220.367
R5180 AVDD.n349 AVDD.t163 220.367
R5181 AVDD.n348 AVDD.t171 220.367
R5182 AVDD.n372 AVDD.t316 220.367
R5183 AVDD.n370 AVDD.t232 220.367
R5184 AVDD.n2892 AVDD.t245 220.367
R5185 AVDD.n2891 AVDD.t142 220.367
R5186 AVDD.n2868 AVDD.t368 220.367
R5187 AVDD.n434 AVDD.t282 220.367
R5188 AVDD.n462 AVDD.t354 220.367
R5189 AVDD.n461 AVDD.t269 220.367
R5190 AVDD.n944 AVDD.t203 220.367
R5191 AVDD.n788 AVDD.t202 220.367
R5192 AVDD.n922 AVDD.t302 220.367
R5193 AVDD.n802 AVDD.t301 220.367
R5194 AVDD.n814 AVDD.t348 220.367
R5195 AVDD.n813 AVDD.t347 220.367
R5196 AVDD.n828 AVDD.t132 220.367
R5197 AVDD.n827 AVDD.t131 220.367
R5198 AVDD.n874 AVDD.t262 220.367
R5199 AVDD.n835 AVDD.t261 220.367
R5200 AVDD.n852 AVDD.t395 220.367
R5201 AVDD.n849 AVDD.t394 220.367
R5202 AVDD.n3290 AVDD.t228 220.367
R5203 AVDD.n104 AVDD.t236 220.367
R5204 AVDD.n119 AVDD.t409 220.367
R5205 AVDD.n117 AVDD.t416 220.367
R5206 AVDD.n3225 AVDD.t267 220.367
R5207 AVDD.n134 AVDD.t277 220.367
R5208 AVDD.n3197 AVDD.t341 220.367
R5209 AVDD.n152 AVDD.t345 220.367
R5210 AVDD.n3155 AVDD.t206 220.367
R5211 AVDD.n3154 AVDD.t210 220.367
R5212 AVDD.n3127 AVDD.t365 220.367
R5213 AVDD.n183 AVDD.t381 220.367
R5214 AVDD.n1342 AVDD.t400 220.367
R5215 AVDD.n1340 AVDD.t404 220.367
R5216 AVDD.n1383 AVDD.t242 220.367
R5217 AVDD.n1325 AVDD.t252 220.367
R5218 AVDD.n1685 AVDD.t374 220.367
R5219 AVDD.n1684 AVDD.t387 220.367
R5220 AVDD.n1408 AVDD.t220 220.367
R5221 AVDD.n1406 AVDD.t230 220.367
R5222 AVDD.n1630 AVDD.t194 220.367
R5223 AVDD.n1629 AVDD.t271 220.367
R5224 AVDD.n1458 AVDD.t313 220.367
R5225 AVDD.n1457 AVDD.t402 220.367
R5226 AVDD.n1563 AVDD.t377 220.367
R5227 AVDD.n1562 AVDD.t392 220.367
R5228 AVDD.n1513 AVDD.t319 220.367
R5229 AVDD.n1511 AVDD.t234 220.367
R5230 AVDD.n2250 AVDD.t248 220.367
R5231 AVDD.n2249 AVDD.t145 220.367
R5232 AVDD.n2285 AVDD.t371 220.367
R5233 AVDD.n2283 AVDD.t286 220.367
R5234 AVDD.n2333 AVDD.t357 220.367
R5235 AVDD.n2217 AVDD.t275 220.367
R5236 AVDD.n1262 AVDD.n1261 204.142
R5237 AVDD.n1287 AVDD.n1286 204.142
R5238 AVDD.n1478 AVDD.n1477 204.142
R5239 AVDD.n388 AVDD.n387 204.142
R5240 AVDD.n2536 AVDD.n2362 204.138
R5241 AVDD.n1262 AVDD.n1260 204.138
R5242 AVDD.n1287 AVDD.n1285 204.138
R5243 AVDD.n1246 AVDD.n1244 204.138
R5244 AVDD.n1478 AVDD.n1476 204.138
R5245 AVDD.n388 AVDD.n386 204.138
R5246 AVDD.n1246 AVDD.n1245 203.763
R5247 AVDD.n1424 AVDD.n1423 203.762
R5248 AVDD.n1313 AVDD.n1312 203.752
R5249 AVDD.n1313 AVDD.n1311 203.381
R5250 AVDD.n1424 AVDD.n1422 203.377
R5251 AVDD.n2605 AVDD.n2604 203.079
R5252 AVDD.n2603 AVDD.n2602 203.079
R5253 AVDD.n2580 AVDD.n2579 203.079
R5254 AVDD.n2539 AVDD.n2538 203.079
R5255 AVDD.n2537 AVDD.n2536 203.079
R5256 AVDD.n2477 AVDD.n2476 203.079
R5257 AVDD.n2475 AVDD.n2472 203.079
R5258 AVDD.n2474 AVDD.n2455 203.079
R5259 AVDD.n2428 AVDD.n2427 203.079
R5260 AVDD.n2426 AVDD.n2425 203.079
R5261 AVDD.n2386 AVDD.n2383 203.079
R5262 AVDD.n1070 AVDD.n1069 203.079
R5263 AVDD.n1068 AVDD.n1067 203.079
R5264 AVDD.n1009 AVDD.n725 203.079
R5265 AVDD.n1011 AVDD.n1010 203.079
R5266 AVDD.n2672 AVDD.n2140 203.079
R5267 AVDD.n2139 AVDD.n2121 203.079
R5268 AVDD.n2138 AVDD.n2104 203.079
R5269 AVDD.n2723 AVDD.n2071 203.079
R5270 AVDD.n2070 AVDD.n2048 203.079
R5271 AVDD.n2069 AVDD.n2034 203.079
R5272 AVDD.n2068 AVDD.n2067 203.079
R5273 AVDD.n2065 AVDD.n2018 203.079
R5274 AVDD.n1975 AVDD.n1974 203.079
R5275 AVDD.n1973 AVDD.n1972 203.079
R5276 AVDD.n1970 AVDD.n1954 203.079
R5277 AVDD.n1883 AVDD.n517 191.802
R5278 AVDD.n537 AVDD.n535 191.802
R5279 AVDD.n1152 AVDD.n1150 191.802
R5280 AVDD.n1178 AVDD.n1176 191.802
R5281 AVDD.n1212 AVDD.n1211 191.802
R5282 AVDD.n1235 AVDD.n1234 191.802
R5283 AVDD.n206 AVDD.n205 191.802
R5284 AVDD.n229 AVDD.n227 191.802
R5285 AVDD.n3051 AVDD.n249 191.802
R5286 AVDD.n269 AVDD.n267 191.802
R5287 AVDD.n3006 AVDD.n289 191.802
R5288 AVDD.n311 AVDD.n309 191.802
R5289 AVDD.n347 AVDD.n346 191.802
R5290 AVDD.n369 AVDD.n368 191.802
R5291 AVDD.n2890 AVDD.n412 191.802
R5292 AVDD.n433 AVDD.n431 191.802
R5293 AVDD.n460 AVDD.n459 191.802
R5294 AVDD.n103 AVDD.n101 191.802
R5295 AVDD.n116 AVDD.n115 191.802
R5296 AVDD.n133 AVDD.n131 191.802
R5297 AVDD.n151 AVDD.n149 191.802
R5298 AVDD.n3153 AVDD.n169 191.802
R5299 AVDD.n182 AVDD.n180 191.802
R5300 AVDD.n1339 AVDD.n1337 191.802
R5301 AVDD.n1324 AVDD.n1323 191.802
R5302 AVDD.n1683 AVDD.n1395 191.802
R5303 AVDD.n1405 AVDD.n1404 191.802
R5304 AVDD.n1628 AVDD.n1441 191.802
R5305 AVDD.n1456 AVDD.n1455 191.802
R5306 AVDD.n1561 AVDD.n1496 191.802
R5307 AVDD.n1510 AVDD.n1509 191.802
R5308 AVDD.n2248 AVDD.n2247 191.802
R5309 AVDD.n2282 AVDD.n2280 191.802
R5310 AVDD.n2216 AVDD.n2214 191.802
R5311 AVDD.n3295 AVDD.n3294 185
R5312 AVDD.n99 AVDD.n96 185
R5313 AVDD.n107 AVDD.n95 185
R5314 AVDD.n3297 AVDD.n95 185
R5315 AVDD.n3286 AVDD.n3285 185
R5316 AVDD.n3278 AVDD.n108 185
R5317 AVDD.n3280 AVDD.n3279 185
R5318 AVDD.n3276 AVDD.n3275 185
R5319 AVDD.n3274 AVDD.n3273 185
R5320 AVDD.n3265 AVDD.n110 185
R5321 AVDD.n3267 AVDD.n3266 185
R5322 AVDD.n3263 AVDD.n3262 185
R5323 AVDD.n3261 AVDD.n3260 185
R5324 AVDD.n3253 AVDD.n113 185
R5325 AVDD.n3255 AVDD.n3254 185
R5326 AVDD.n3251 AVDD.n3250 185
R5327 AVDD.n3249 AVDD.n3248 185
R5328 AVDD.n3241 AVDD.n123 185
R5329 AVDD.n3243 AVDD.n3242 185
R5330 AVDD.n3234 AVDD.n126 185
R5331 AVDD.n3236 AVDD.n3235 185
R5332 AVDD.n3232 AVDD.n3231 185
R5333 AVDD.n3230 AVDD.n3229 185
R5334 AVDD.n137 AVDD.n129 185
R5335 AVDD.n139 AVDD.n138 185
R5336 AVDD.n3221 AVDD.n3220 185
R5337 AVDD.n3219 AVDD.n3218 185
R5338 AVDD.n3216 AVDD.n3215 185
R5339 AVDD.n3214 AVDD.n3213 185
R5340 AVDD.n3206 AVDD.n141 185
R5341 AVDD.n3208 AVDD.n3207 185
R5342 AVDD.n3204 AVDD.n3203 185
R5343 AVDD.n3202 AVDD.n3201 185
R5344 AVDD.n155 AVDD.n146 185
R5345 AVDD.n157 AVDD.n156 185
R5346 AVDD.n3193 AVDD.n3192 185
R5347 AVDD.n3191 AVDD.n3190 185
R5348 AVDD.n3183 AVDD.n159 185
R5349 AVDD.n3185 AVDD.n3184 185
R5350 AVDD.n3181 AVDD.n3180 185
R5351 AVDD.n3179 AVDD.n3178 185
R5352 AVDD.n3171 AVDD.n162 185
R5353 AVDD.n3173 AVDD.n3172 185
R5354 AVDD.n3169 AVDD.n3168 185
R5355 AVDD.n3167 AVDD.n3166 185
R5356 AVDD.n3159 AVDD.n166 185
R5357 AVDD.n3161 AVDD.n3160 185
R5358 AVDD.n3148 AVDD.n168 185
R5359 AVDD.n3150 AVDD.n3149 185
R5360 AVDD.n3146 AVDD.n3145 185
R5361 AVDD.n3144 AVDD.n3143 185
R5362 AVDD.n3136 AVDD.n172 185
R5363 AVDD.n3138 AVDD.n3137 185
R5364 AVDD.n3134 AVDD.n3133 185
R5365 AVDD.n3132 AVDD.n3131 185
R5366 AVDD.n3121 AVDD.n177 185
R5367 AVDD.n3123 AVDD.n3122 185
R5368 AVDD.n3119 AVDD.n3118 185
R5369 AVDD.n3117 AVDD.n3116 185
R5370 AVDD.n188 AVDD.n187 185
R5371 AVDD.n3110 AVDD.n42 185
R5372 AVDD.n3297 AVDD.n42 185
R5373 AVDD.n192 AVDD.n94 185
R5374 AVDD.n3297 AVDD.n94 185
R5375 AVDD.n1334 AVDD.n1333 185
R5376 AVDD.n1347 AVDD.n1346 185
R5377 AVDD.n1349 AVDD.n1348 185
R5378 AVDD.n1353 AVDD.n1352 185
R5379 AVDD.n1351 AVDD.n1330 185
R5380 AVDD.n1360 AVDD.n1359 185
R5381 AVDD.n1362 AVDD.n1361 185
R5382 AVDD.n1366 AVDD.n1365 185
R5383 AVDD.n1364 AVDD.n1328 185
R5384 AVDD.n1373 AVDD.n1372 185
R5385 AVDD.n1375 AVDD.n1374 185
R5386 AVDD.n1379 AVDD.n1378 185
R5387 AVDD.n1377 AVDD.n1321 185
R5388 AVDD.n1388 AVDD.n1387 185
R5389 AVDD.n1390 AVDD.n1389 185
R5390 AVDD.n1699 AVDD.n1698 185
R5391 AVDD.n1697 AVDD.n1696 185
R5392 AVDD.n1689 AVDD.n1392 185
R5393 AVDD.n1691 AVDD.n1690 185
R5394 AVDD.n1678 AVDD.n1394 185
R5395 AVDD.n1680 AVDD.n1679 185
R5396 AVDD.n1671 AVDD.n1397 185
R5397 AVDD.n1673 AVDD.n1672 185
R5398 AVDD.n1669 AVDD.n1668 185
R5399 AVDD.n1667 AVDD.n1666 185
R5400 AVDD.n1658 AVDD.n1399 185
R5401 AVDD.n1660 AVDD.n1659 185
R5402 AVDD.n1656 AVDD.n1655 185
R5403 AVDD.n1654 AVDD.n1653 185
R5404 AVDD.n1646 AVDD.n1402 185
R5405 AVDD.n1648 AVDD.n1647 185
R5406 AVDD.n1639 AVDD.n1435 185
R5407 AVDD.n1641 AVDD.n1640 185
R5408 AVDD.n1637 AVDD.n1636 185
R5409 AVDD.n1635 AVDD.n1634 185
R5410 AVDD.n1623 AVDD.n1438 185
R5411 AVDD.n1625 AVDD.n1624 185
R5412 AVDD.n1444 AVDD.n1443 185
R5413 AVDD.n1618 AVDD.n62 185
R5414 AVDD.n3297 AVDD.n62 185
R5415 AVDD.n1446 AVDD.n93 185
R5416 AVDD.n3297 AVDD.n93 185
R5417 AVDD.n1614 AVDD.n1613 185
R5418 AVDD.n1449 AVDD.n1447 185
R5419 AVDD.n1451 AVDD.n1450 185
R5420 AVDD.n1608 AVDD.n1607 185
R5421 AVDD.n1606 AVDD.n1605 185
R5422 AVDD.n1598 AVDD.n1453 185
R5423 AVDD.n1600 AVDD.n1599 185
R5424 AVDD.n1596 AVDD.n1595 185
R5425 AVDD.n1594 AVDD.n1593 185
R5426 AVDD.n1586 AVDD.n1462 185
R5427 AVDD.n1588 AVDD.n1587 185
R5428 AVDD.n1579 AVDD.n1489 185
R5429 AVDD.n1581 AVDD.n1580 185
R5430 AVDD.n1577 AVDD.n1576 185
R5431 AVDD.n1575 AVDD.n1574 185
R5432 AVDD.n1567 AVDD.n1492 185
R5433 AVDD.n1569 AVDD.n1568 185
R5434 AVDD.n1556 AVDD.n1495 185
R5435 AVDD.n1558 AVDD.n1557 185
R5436 AVDD.n1500 AVDD.n1498 185
R5437 AVDD.n1502 AVDD.n1501 185
R5438 AVDD.n1551 AVDD.n1550 185
R5439 AVDD.n1549 AVDD.n1548 185
R5440 AVDD.n1540 AVDD.n1504 185
R5441 AVDD.n1542 AVDD.n1541 185
R5442 AVDD.n1538 AVDD.n1537 185
R5443 AVDD.n1536 AVDD.n1535 185
R5444 AVDD.n1528 AVDD.n1507 185
R5445 AVDD.n1530 AVDD.n1529 185
R5446 AVDD.n1526 AVDD.n1525 185
R5447 AVDD.n1524 AVDD.n1523 185
R5448 AVDD.n1519 AVDD.n1518 185
R5449 AVDD.n12 AVDD.n9 185
R5450 AVDD.n3300 AVDD.n3299 185
R5451 AVDD.n2235 AVDD.n11 185
R5452 AVDD.n2239 AVDD.n2238 185
R5453 AVDD.n2241 AVDD.n2240 185
R5454 AVDD.n2244 AVDD.n2243 185
R5455 AVDD.n2242 AVDD.n2232 185
R5456 AVDD.n2256 AVDD.n2255 185
R5457 AVDD.n2254 AVDD.n2230 185
R5458 AVDD.n2264 AVDD.n2263 185
R5459 AVDD.n2266 AVDD.n2265 185
R5460 AVDD.n2270 AVDD.n2269 185
R5461 AVDD.n2268 AVDD.n2227 185
R5462 AVDD.n2277 AVDD.n2276 185
R5463 AVDD.n2275 AVDD.n2225 185
R5464 AVDD.n2290 AVDD.n2289 185
R5465 AVDD.n2292 AVDD.n2291 185
R5466 AVDD.n2296 AVDD.n2295 185
R5467 AVDD.n2294 AVDD.n2222 185
R5468 AVDD.n2303 AVDD.n2302 185
R5469 AVDD.n2305 AVDD.n2304 185
R5470 AVDD.n2309 AVDD.n2308 185
R5471 AVDD.n2307 AVDD.n2219 185
R5472 AVDD.n2315 AVDD.n2314 185
R5473 AVDD.n2317 AVDD.n2316 185
R5474 AVDD.n2327 AVDD.n2319 185
R5475 AVDD.n2329 AVDD.n2328 185
R5476 AVDD.n2325 AVDD.n2324 185
R5477 AVDD.n2322 AVDD.n92 185
R5478 AVDD.n3297 AVDD.n92 185
R5479 AVDD.n2187 AVDD.n2185 185
R5480 AVDD.n2185 AVDD.n13 185
R5481 AVDD.n2640 AVDD.n2639 185
R5482 AVDD.n2643 AVDD.n2640 185
R5483 AVDD.n2193 AVDD.n2184 185
R5484 AVDD.n2644 AVDD.n2184 185
R5485 AVDD.n2192 AVDD.n2183 185
R5486 AVDD.n2645 AVDD.n2183 185
R5487 AVDD.n2199 AVDD.n2198 185
R5488 AVDD.n2199 AVDD.n2182 185
R5489 AVDD.n2201 AVDD.n2200 185
R5490 AVDD.n2202 AVDD.n2201 185
R5491 AVDD.n2209 AVDD.n2208 185
R5492 AVDD.n2208 AVDD.n2207 185
R5493 AVDD.n2197 AVDD.n2196 185
R5494 AVDD.n2197 AVDD.n2165 185
R5495 AVDD.n2635 AVDD.n2164 185
R5496 AVDD.n2653 AVDD.n2164 185
R5497 AVDD.n2634 AVDD.n2163 185
R5498 AVDD.n2654 AVDD.n2163 185
R5499 AVDD.n2211 AVDD.n2162 185
R5500 AVDD.n2655 AVDD.n2162 185
R5501 AVDD.n2624 AVDD.n2623 185
R5502 AVDD.n2623 AVDD.n2161 185
R5503 AVDD.n2622 AVDD.n2621 185
R5504 AVDD.n2622 AVDD.n2147 185
R5505 AVDD.n2338 AVDD.n2146 185
R5506 AVDD.n2665 AVDD.n2146 185
R5507 AVDD.n2613 AVDD.n2145 185
R5508 AVDD.n2666 AVDD.n2145 185
R5509 AVDD.n2611 AVDD.n2144 185
R5510 AVDD.n2667 AVDD.n2144 185
R5511 AVDD.n2609 AVDD.n2608 185
R5512 AVDD.n2608 AVDD.n2128 185
R5513 AVDD.n2341 AVDD.n2127 185
R5514 AVDD.n2677 AVDD.n2127 185
R5515 AVDD.n2599 AVDD.n2126 185
R5516 AVDD.n2678 AVDD.n2126 185
R5517 AVDD.n2596 AVDD.n2125 185
R5518 AVDD.n2679 AVDD.n2125 185
R5519 AVDD.n2594 AVDD.n2593 185
R5520 AVDD.n2593 AVDD.n2124 185
R5521 AVDD.n2346 AVDD.n2113 185
R5522 AVDD.n2690 AVDD.n2113 185
R5523 AVDD.n2585 AVDD.n2112 185
R5524 AVDD.n2691 AVDD.n2112 185
R5525 AVDD.n2583 AVDD.n2111 185
R5526 AVDD.n2692 AVDD.n2111 185
R5527 AVDD.n2567 AVDD.n2348 185
R5528 AVDD.n2567 AVDD.n2110 185
R5529 AVDD.n2569 AVDD.n2568 185
R5530 AVDD.n2568 AVDD.n2096 185
R5531 AVDD.n2565 AVDD.n2095 185
R5532 AVDD.n2704 AVDD.n2095 185
R5533 AVDD.n2563 AVDD.n2094 185
R5534 AVDD.n2705 AVDD.n2094 185
R5535 AVDD.n2355 AVDD.n2093 185
R5536 AVDD.n2706 AVDD.n2093 185
R5537 AVDD.n2558 AVDD.n2557 185
R5538 AVDD.n2557 AVDD.n2092 185
R5539 AVDD.n2556 AVDD.n2555 185
R5540 AVDD.n2556 AVDD.n2078 185
R5541 AVDD.n2357 AVDD.n2077 185
R5542 AVDD.n2716 AVDD.n2077 185
R5543 AVDD.n2547 AVDD.n2076 185
R5544 AVDD.n2717 AVDD.n2076 185
R5545 AVDD.n2545 AVDD.n2075 185
R5546 AVDD.n2718 AVDD.n2075 185
R5547 AVDD.n2543 AVDD.n2542 185
R5548 AVDD.n2542 AVDD.n2055 185
R5549 AVDD.n2360 AVDD.n2054 185
R5550 AVDD.n2728 AVDD.n2054 185
R5551 AVDD.n2533 AVDD.n2053 185
R5552 AVDD.n2729 AVDD.n2053 185
R5553 AVDD.n2528 AVDD.n2052 185
R5554 AVDD.n2730 AVDD.n2052 185
R5555 AVDD.n2366 AVDD.n2365 185
R5556 AVDD.n2365 AVDD.n2051 185
R5557 AVDD.n2486 AVDD.n2040 185
R5558 AVDD.n2741 AVDD.n2040 185
R5559 AVDD.n2481 AVDD.n2039 185
R5560 AVDD.n2742 AVDD.n2039 185
R5561 AVDD.n2491 AVDD.n2038 185
R5562 AVDD.n2743 AVDD.n2038 185
R5563 AVDD.n2480 AVDD.n2479 185
R5564 AVDD.n2479 AVDD.n2037 185
R5565 AVDD.n2471 AVDD.n2028 185
R5566 AVDD.n2754 AVDD.n2028 185
R5567 AVDD.n2499 AVDD.n2027 185
R5568 AVDD.n2755 AVDD.n2027 185
R5569 AVDD.n2501 AVDD.n2026 185
R5570 AVDD.n2756 AVDD.n2026 185
R5571 AVDD.n2470 AVDD.n2469 185
R5572 AVDD.n2469 AVDD.n2025 185
R5573 AVDD.n2468 AVDD.n2463 185
R5574 AVDD.n2468 AVDD.n2467 185
R5575 AVDD.n2462 AVDD.n2458 185
R5576 AVDD.n2462 AVDD.n2009 185
R5577 AVDD.n2509 AVDD.n2008 185
R5578 AVDD.n2768 AVDD.n2008 185
R5579 AVDD.n2457 AVDD.n2007 185
R5580 AVDD.n2769 AVDD.n2007 185
R5581 AVDD.n2453 AVDD.n2006 185
R5582 AVDD.n2770 AVDD.n2006 185
R5583 AVDD.n2518 AVDD.n2517 185
R5584 AVDD.n2517 AVDD.n1996 185
R5585 AVDD.n2452 AVDD.n1995 185
R5586 AVDD.n2780 AVDD.n1995 185
R5587 AVDD.n2450 AVDD.n1994 185
R5588 AVDD.n2781 AVDD.n1994 185
R5589 AVDD.n2371 AVDD.n1993 185
R5590 AVDD.n2782 AVDD.n1993 185
R5591 AVDD.n2441 AVDD.n2440 185
R5592 AVDD.n2440 AVDD.n1981 185
R5593 AVDD.n2373 AVDD.n1982 185
R5594 AVDD.t16 AVDD.n1982 185
R5595 AVDD.n2433 AVDD.n1980 185
R5596 AVDD.n2793 AVDD.n1980 185
R5597 AVDD.n2431 AVDD.n1979 185
R5598 AVDD.n2794 AVDD.n1979 185
R5599 AVDD.n2376 AVDD.n2375 185
R5600 AVDD.n2375 AVDD.n1978 185
R5601 AVDD.n2422 AVDD.n1964 185
R5602 AVDD.n2805 AVDD.n1964 185
R5603 AVDD.n2419 AVDD.n1963 185
R5604 AVDD.n2806 AVDD.n1963 185
R5605 AVDD.n2417 AVDD.n1962 185
R5606 AVDD.n2807 AVDD.n1962 185
R5607 AVDD.n2402 AVDD.n2381 185
R5608 AVDD.n2402 AVDD.n1961 185
R5609 AVDD.n2407 AVDD.n2401 185
R5610 AVDD.n2407 AVDD.n2406 185
R5611 AVDD.n2409 AVDD.n2408 185
R5612 AVDD.n2408 AVDD.n1945 185
R5613 AVDD.n2399 AVDD.n1944 185
R5614 AVDD.n2819 AVDD.n1944 185
R5615 AVDD.n2384 AVDD.n1943 185
R5616 AVDD.n2820 AVDD.n1943 185
R5617 AVDD.n2391 AVDD.n1942 185
R5618 AVDD.n2821 AVDD.n1942 185
R5619 AVDD.n2389 AVDD.n470 185
R5620 AVDD.n472 AVDD.n470 185
R5621 AVDD.n2832 AVDD.n2831 185
R5622 AVDD.n2831 AVDD.n2830 185
R5623 AVDD.n469 AVDD.n467 185
R5624 AVDD.n471 AVDD.n469 185
R5625 AVDD.n1930 AVDD.n1929 185
R5626 AVDD.n1931 AVDD.n1930 185
R5627 AVDD.n482 AVDD.n481 185
R5628 AVDD.n481 AVDD.n480 185
R5629 AVDD.n1913 AVDD.n1912 185
R5630 AVDD.n1914 AVDD.n1913 185
R5631 AVDD.n1911 AVDD.n1901 185
R5632 AVDD.n1911 AVDD.n1910 185
R5633 AVDD.n1900 AVDD.n1899 185
R5634 AVDD.n1909 AVDD.n1900 185
R5635 AVDD.n1903 AVDD.n1902 185
R5636 AVDD.n1904 AVDD.n1903 185
R5637 AVDD.n500 AVDD.n499 185
R5638 AVDD.n502 AVDD.n500 185
R5639 AVDD.n1924 AVDD.n1923 185
R5640 AVDD.n1923 AVDD.n1922 185
R5641 AVDD.n498 AVDD.n490 185
R5642 AVDD.n501 AVDD.n498 185
R5643 AVDD.n497 AVDD.n496 185
R5644 AVDD.n457 AVDD.n456 185
R5645 AVDD.n2842 AVDD.n2841 185
R5646 AVDD.n2845 AVDD.n2844 185
R5647 AVDD.n455 AVDD.n452 185
R5648 AVDD.n449 AVDD.n447 185
R5649 AVDD.n2851 AVDD.n2850 185
R5650 AVDD.n2853 AVDD.n446 185
R5651 AVDD.n2855 AVDD.n2854 185
R5652 AVDD.n442 AVDD.n441 185
R5653 AVDD.n2861 AVDD.n2860 185
R5654 AVDD.n2864 AVDD.n2863 185
R5655 AVDD.n440 AVDD.n437 185
R5656 AVDD.n428 AVDD.n426 185
R5657 AVDD.n2873 AVDD.n2872 185
R5658 AVDD.n2875 AVDD.n425 185
R5659 AVDD.n2877 AVDD.n2876 185
R5660 AVDD.n419 AVDD.n417 185
R5661 AVDD.n2883 AVDD.n2882 185
R5662 AVDD.n2885 AVDD.n416 185
R5663 AVDD.n2887 AVDD.n2886 185
R5664 AVDD.n410 AVDD.n409 185
R5665 AVDD.n2897 AVDD.n2896 185
R5666 AVDD.n2899 AVDD.n408 185
R5667 AVDD.n2901 AVDD.n2900 185
R5668 AVDD.n402 AVDD.n400 185
R5669 AVDD.n2907 AVDD.n2906 185
R5670 AVDD.n2909 AVDD.n399 185
R5671 AVDD.n2911 AVDD.n2910 185
R5672 AVDD.n380 AVDD.n378 185
R5673 AVDD.n2917 AVDD.n2916 185
R5674 AVDD.n2919 AVDD.n377 185
R5675 AVDD.n2921 AVDD.n2920 185
R5676 AVDD.n366 AVDD.n364 185
R5677 AVDD.n2927 AVDD.n2926 185
R5678 AVDD.n2929 AVDD.n363 185
R5679 AVDD.n2931 AVDD.n2930 185
R5680 AVDD.n359 AVDD.n358 185
R5681 AVDD.n2938 AVDD.n2937 185
R5682 AVDD.n2941 AVDD.n2940 185
R5683 AVDD.n357 AVDD.n354 185
R5684 AVDD.n344 AVDD.n342 185
R5685 AVDD.n2947 AVDD.n2946 185
R5686 AVDD.n2949 AVDD.n341 185
R5687 AVDD.n2951 AVDD.n2950 185
R5688 AVDD.n336 AVDD.n334 185
R5689 AVDD.n2957 AVDD.n2956 185
R5690 AVDD.n2959 AVDD.n333 185
R5691 AVDD.n2961 AVDD.n2960 185
R5692 AVDD.n327 AVDD.n325 185
R5693 AVDD.n2967 AVDD.n2966 185
R5694 AVDD.n2969 AVDD.n324 185
R5695 AVDD.n2971 AVDD.n2970 185
R5696 AVDD.n320 AVDD.n319 185
R5697 AVDD.n2977 AVDD.n2976 185
R5698 AVDD.n2980 AVDD.n2979 185
R5699 AVDD.n318 AVDD.n315 185
R5700 AVDD.n307 AVDD.n306 185
R5701 AVDD.n2989 AVDD.n2988 185
R5702 AVDD.n2991 AVDD.n305 185
R5703 AVDD.n2993 AVDD.n2992 185
R5704 AVDD.n303 AVDD.n297 185
R5705 AVDD.n2999 AVDD.n2998 185
R5706 AVDD.n3001 AVDD.n293 185
R5707 AVDD.n3003 AVDD.n3002 185
R5708 AVDD.n286 AVDD.n284 185
R5709 AVDD.n3013 AVDD.n3012 185
R5710 AVDD.n3015 AVDD.n283 185
R5711 AVDD.n3017 AVDD.n3016 185
R5712 AVDD.n278 AVDD.n277 185
R5713 AVDD.n3023 AVDD.n3022 185
R5714 AVDD.n3026 AVDD.n3025 185
R5715 AVDD.n276 AVDD.n273 185
R5716 AVDD.n265 AVDD.n264 185
R5717 AVDD.n3035 AVDD.n3034 185
R5718 AVDD.n3038 AVDD.n3037 185
R5719 AVDD.n263 AVDD.n260 185
R5720 AVDD.n256 AVDD.n254 185
R5721 AVDD.n3044 AVDD.n3043 185
R5722 AVDD.n3046 AVDD.n253 185
R5723 AVDD.n3048 AVDD.n3047 185
R5724 AVDD.n246 AVDD.n244 185
R5725 AVDD.n3058 AVDD.n3057 185
R5726 AVDD.n3060 AVDD.n243 185
R5727 AVDD.n3062 AVDD.n3061 185
R5728 AVDD.n238 AVDD.n237 185
R5729 AVDD.n3068 AVDD.n3067 185
R5730 AVDD.n3071 AVDD.n3070 185
R5731 AVDD.n236 AVDD.n233 185
R5732 AVDD.n224 AVDD.n222 185
R5733 AVDD.n3080 AVDD.n3079 185
R5734 AVDD.n3082 AVDD.n221 185
R5735 AVDD.n3084 AVDD.n3083 185
R5736 AVDD.n216 AVDD.n215 185
R5737 AVDD.n3090 AVDD.n3089 185
R5738 AVDD.n3092 AVDD.n214 185
R5739 AVDD.n3094 AVDD.n3093 185
R5740 AVDD.n203 AVDD.n201 185
R5741 AVDD.n3100 AVDD.n3099 185
R5742 AVDD.n3102 AVDD.n199 185
R5743 AVDD.n3104 AVDD.n3103 185
R5744 AVDD.n1732 AVDD.n193 185
R5745 AVDD.n1735 AVDD.n194 185
R5746 AVDD.n1737 AVDD.n1731 185
R5747 AVDD.n1739 AVDD.n1738 185
R5748 AVDD.n1231 AVDD.n1229 185
R5749 AVDD.n1745 AVDD.n1744 185
R5750 AVDD.n1747 AVDD.n1228 185
R5751 AVDD.n1749 AVDD.n1748 185
R5752 AVDD.n1223 AVDD.n1221 185
R5753 AVDD.n1756 AVDD.n1755 185
R5754 AVDD.n1758 AVDD.n1220 185
R5755 AVDD.n1760 AVDD.n1759 185
R5756 AVDD.n1209 AVDD.n1207 185
R5757 AVDD.n1767 AVDD.n1766 185
R5758 AVDD.n1769 AVDD.n1206 185
R5759 AVDD.n1771 AVDD.n1770 185
R5760 AVDD.n1202 AVDD.n1201 185
R5761 AVDD.n1777 AVDD.n1776 185
R5762 AVDD.n1779 AVDD.n1200 185
R5763 AVDD.n1781 AVDD.n1780 185
R5764 AVDD.n1194 AVDD.n1192 185
R5765 AVDD.n1787 AVDD.n1786 185
R5766 AVDD.n1789 AVDD.n1191 185
R5767 AVDD.n1791 AVDD.n1790 185
R5768 AVDD.n1187 AVDD.n1186 185
R5769 AVDD.n1797 AVDD.n1796 185
R5770 AVDD.n1800 AVDD.n1799 185
R5771 AVDD.n1185 AVDD.n1182 185
R5772 AVDD.n1173 AVDD.n1171 185
R5773 AVDD.n1809 AVDD.n1808 185
R5774 AVDD.n1811 AVDD.n1170 185
R5775 AVDD.n1813 AVDD.n1812 185
R5776 AVDD.n1164 AVDD.n1162 185
R5777 AVDD.n1819 AVDD.n1818 185
R5778 AVDD.n1821 AVDD.n1161 185
R5779 AVDD.n1822 AVDD.n1157 185
R5780 AVDD.n1825 AVDD.n1824 185
R5781 AVDD.n1159 AVDD.n1156 185
R5782 AVDD.n1148 AVDD.n1146 185
R5783 AVDD.n1834 AVDD.n1833 185
R5784 AVDD.n1836 AVDD.n1145 185
R5785 AVDD.n1838 AVDD.n1837 185
R5786 AVDD.n553 AVDD.n551 185
R5787 AVDD.n1845 AVDD.n1844 185
R5788 AVDD.n1847 AVDD.n550 185
R5789 AVDD.n1849 AVDD.n1848 185
R5790 AVDD.n546 AVDD.n545 185
R5791 AVDD.n1855 AVDD.n1854 185
R5792 AVDD.n1858 AVDD.n1857 185
R5793 AVDD.n544 AVDD.n541 185
R5794 AVDD.n533 AVDD.n532 185
R5795 AVDD.n1867 AVDD.n1866 185
R5796 AVDD.n1870 AVDD.n1869 185
R5797 AVDD.n531 AVDD.n528 185
R5798 AVDD.n524 AVDD.n522 185
R5799 AVDD.n1876 AVDD.n1875 185
R5800 AVDD.n1878 AVDD.n521 185
R5801 AVDD.n1880 AVDD.n1879 185
R5802 AVDD.n514 AVDD.n513 185
R5803 AVDD.n1890 AVDD.n1889 185
R5804 AVDD.n1893 AVDD.n1892 185
R5805 AVDD.n511 AVDD.n503 185
R5806 AVDD.n503 AVDD.n501 185
R5807 AVDD.n1921 AVDD.n1920 185
R5808 AVDD.n1922 AVDD.n1921 185
R5809 AVDD.n506 AVDD.n504 185
R5810 AVDD.n504 AVDD.n502 185
R5811 AVDD.n1906 AVDD.n1905 185
R5812 AVDD.n1906 AVDD.n1904 185
R5813 AVDD.n1908 AVDD.n1907 185
R5814 AVDD.n1909 AVDD.n1908 185
R5815 AVDD.n1898 AVDD.n1897 185
R5816 AVDD.n1910 AVDD.n1898 185
R5817 AVDD.n1916 AVDD.n1915 185
R5818 AVDD.n1915 AVDD.n1914 185
R5819 AVDD.n509 AVDD.n479 185
R5820 AVDD.n480 AVDD.n479 185
R5821 AVDD.n1933 AVDD.n1932 185
R5822 AVDD.n1932 AVDD.n1931 185
R5823 AVDD.n1934 AVDD.n473 185
R5824 AVDD.n473 AVDD.n471 185
R5825 AVDD.n2829 AVDD.n2828 185
R5826 AVDD.n2830 AVDD.n2829 185
R5827 AVDD.n476 AVDD.n474 185
R5828 AVDD.n474 AVDD.n472 185
R5829 AVDD.n2823 AVDD.n2822 185
R5830 AVDD.n2822 AVDD.n2821 185
R5831 AVDD.n1947 AVDD.n1941 185
R5832 AVDD.n2820 AVDD.n1941 185
R5833 AVDD.n2818 AVDD.n2817 185
R5834 AVDD.n2819 AVDD.n2818 185
R5835 AVDD.n1949 AVDD.n1946 185
R5836 AVDD.n1946 AVDD.n1945 185
R5837 AVDD.n2405 AVDD.n2404 185
R5838 AVDD.n2406 AVDD.n2405 185
R5839 AVDD.n1959 AVDD.n1957 185
R5840 AVDD.n1961 AVDD.n1959 185
R5841 AVDD.n2809 AVDD.n2808 185
R5842 AVDD.n2808 AVDD.n2807 185
R5843 AVDD.n1966 AVDD.n1960 185
R5844 AVDD.n2806 AVDD.n1960 185
R5845 AVDD.n2804 AVDD.n2803 185
R5846 AVDD.n2805 AVDD.n2804 185
R5847 AVDD.n1968 AVDD.n1965 185
R5848 AVDD.n1978 AVDD.n1965 185
R5849 AVDD.n2796 AVDD.n2795 185
R5850 AVDD.n2795 AVDD.n2794 185
R5851 AVDD.n1984 AVDD.n1977 185
R5852 AVDD.n2793 AVDD.n1977 185
R5853 AVDD.n2792 AVDD.n2791 185
R5854 AVDD.t16 AVDD.n2792 185
R5855 AVDD.n1986 AVDD.n1983 185
R5856 AVDD.n1983 AVDD.n1981 185
R5857 AVDD.n2784 AVDD.n2783 185
R5858 AVDD.n2783 AVDD.n2782 185
R5859 AVDD.n1998 AVDD.n1992 185
R5860 AVDD.n2781 AVDD.n1992 185
R5861 AVDD.n2779 AVDD.n2778 185
R5862 AVDD.n2780 AVDD.n2779 185
R5863 AVDD.n2000 AVDD.n1997 185
R5864 AVDD.n1997 AVDD.n1996 185
R5865 AVDD.n2772 AVDD.n2771 185
R5866 AVDD.n2771 AVDD.n2770 185
R5867 AVDD.n2011 AVDD.n2005 185
R5868 AVDD.n2769 AVDD.n2005 185
R5869 AVDD.n2767 AVDD.n2766 185
R5870 AVDD.n2768 AVDD.n2767 185
R5871 AVDD.n2013 AVDD.n2010 185
R5872 AVDD.n2010 AVDD.n2009 185
R5873 AVDD.n2466 AVDD.n2465 185
R5874 AVDD.n2467 AVDD.n2466 185
R5875 AVDD.n2023 AVDD.n2021 185
R5876 AVDD.n2025 AVDD.n2023 185
R5877 AVDD.n2758 AVDD.n2757 185
R5878 AVDD.n2757 AVDD.n2756 185
R5879 AVDD.n2030 AVDD.n2024 185
R5880 AVDD.n2755 AVDD.n2024 185
R5881 AVDD.n2753 AVDD.n2752 185
R5882 AVDD.n2754 AVDD.n2753 185
R5883 AVDD.n2032 AVDD.n2029 185
R5884 AVDD.n2037 AVDD.n2029 185
R5885 AVDD.n2745 AVDD.n2744 185
R5886 AVDD.n2744 AVDD.n2743 185
R5887 AVDD.n2042 AVDD.n2036 185
R5888 AVDD.n2742 AVDD.n2036 185
R5889 AVDD.n2740 AVDD.n2739 185
R5890 AVDD.n2741 AVDD.n2740 185
R5891 AVDD.n2044 AVDD.n2041 185
R5892 AVDD.n2051 AVDD.n2041 185
R5893 AVDD.n2732 AVDD.n2731 185
R5894 AVDD.n2731 AVDD.n2730 185
R5895 AVDD.n2057 AVDD.n2050 185
R5896 AVDD.n2729 AVDD.n2050 185
R5897 AVDD.n2727 AVDD.n2726 185
R5898 AVDD.n2728 AVDD.n2727 185
R5899 AVDD.n2059 AVDD.n2056 185
R5900 AVDD.n2056 AVDD.n2055 185
R5901 AVDD.n2720 AVDD.n2719 185
R5902 AVDD.n2719 AVDD.n2718 185
R5903 AVDD.n2080 AVDD.n2074 185
R5904 AVDD.n2717 AVDD.n2074 185
R5905 AVDD.n2715 AVDD.n2714 185
R5906 AVDD.n2716 AVDD.n2715 185
R5907 AVDD.n2082 AVDD.n2079 185
R5908 AVDD.n2079 AVDD.n2078 185
R5909 AVDD.n2090 AVDD.n2088 185
R5910 AVDD.n2092 AVDD.n2090 185
R5911 AVDD.n2708 AVDD.n2707 185
R5912 AVDD.n2707 AVDD.n2706 185
R5913 AVDD.n2098 AVDD.n2091 185
R5914 AVDD.n2705 AVDD.n2091 185
R5915 AVDD.n2703 AVDD.n2702 185
R5916 AVDD.n2704 AVDD.n2703 185
R5917 AVDD.n2100 AVDD.n2097 185
R5918 AVDD.n2097 AVDD.n2096 185
R5919 AVDD.n2108 AVDD.n2106 185
R5920 AVDD.n2110 AVDD.n2108 185
R5921 AVDD.n2694 AVDD.n2693 185
R5922 AVDD.n2693 AVDD.n2692 185
R5923 AVDD.n2115 AVDD.n2109 185
R5924 AVDD.n2691 AVDD.n2109 185
R5925 AVDD.n2689 AVDD.n2688 185
R5926 AVDD.n2690 AVDD.n2689 185
R5927 AVDD.n2117 AVDD.n2114 185
R5928 AVDD.n2124 AVDD.n2114 185
R5929 AVDD.n2681 AVDD.n2680 185
R5930 AVDD.n2680 AVDD.n2679 185
R5931 AVDD.n2130 AVDD.n2123 185
R5932 AVDD.n2678 AVDD.n2123 185
R5933 AVDD.n2676 AVDD.n2675 185
R5934 AVDD.n2677 AVDD.n2676 185
R5935 AVDD.n2132 AVDD.n2129 185
R5936 AVDD.n2129 AVDD.n2128 185
R5937 AVDD.n2669 AVDD.n2668 185
R5938 AVDD.n2668 AVDD.n2667 185
R5939 AVDD.n2149 AVDD.n2143 185
R5940 AVDD.n2666 AVDD.n2143 185
R5941 AVDD.n2664 AVDD.n2663 185
R5942 AVDD.n2665 AVDD.n2664 185
R5943 AVDD.n2151 AVDD.n2148 185
R5944 AVDD.n2148 AVDD.n2147 185
R5945 AVDD.n2159 AVDD.n2157 185
R5946 AVDD.n2161 AVDD.n2159 185
R5947 AVDD.n2657 AVDD.n2656 185
R5948 AVDD.n2656 AVDD.n2655 185
R5949 AVDD.n2167 AVDD.n2160 185
R5950 AVDD.n2654 AVDD.n2160 185
R5951 AVDD.n2652 AVDD.n2651 185
R5952 AVDD.n2653 AVDD.n2652 185
R5953 AVDD.n2169 AVDD.n2166 185
R5954 AVDD.n2166 AVDD.n2165 185
R5955 AVDD.n2206 AVDD.n2205 185
R5956 AVDD.n2207 AVDD.n2206 185
R5957 AVDD.n2204 AVDD.n2203 185
R5958 AVDD.n2204 AVDD.n2202 185
R5959 AVDD.n2179 AVDD.n2178 185
R5960 AVDD.n2182 AVDD.n2179 185
R5961 AVDD.n2647 AVDD.n2646 185
R5962 AVDD.n2646 AVDD.n2645 185
R5963 AVDD.n2181 AVDD.n2180 185
R5964 AVDD.n2644 AVDD.n2181 185
R5965 AVDD.n2642 AVDD.n2641 185
R5966 AVDD.n2643 AVDD.n2642 185
R5967 AVDD.n2175 AVDD.n97 185
R5968 AVDD.n97 AVDD.n13 185
R5969 AVDD.n775 AVDD.n774 185
R5970 AVDD.n847 AVDD.n846 185
R5971 AVDD.n857 AVDD.n856 185
R5972 AVDD.n860 AVDD.n859 185
R5973 AVDD.n844 AVDD.n840 185
R5974 AVDD.n866 AVDD.n865 185
R5975 AVDD.n871 AVDD.n870 185
R5976 AVDD.n868 AVDD.n837 185
R5977 AVDD.n867 AVDD.n833 185
R5978 AVDD.n879 AVDD.n878 185
R5979 AVDD.n882 AVDD.n881 185
R5980 AVDD.n825 AVDD.n824 185
R5981 AVDD.n888 AVDD.n887 185
R5982 AVDD.n891 AVDD.n890 185
R5983 AVDD.n823 AVDD.n819 185
R5984 AVDD.n897 AVDD.n896 185
R5985 AVDD.n900 AVDD.n899 185
R5986 AVDD.n811 AVDD.n810 185
R5987 AVDD.n907 AVDD.n906 185
R5988 AVDD.n910 AVDD.n909 185
R5989 AVDD.n809 AVDD.n806 185
R5990 AVDD.n916 AVDD.n915 185
R5991 AVDD.n919 AVDD.n918 185
R5992 AVDD.n799 AVDD.n797 185
R5993 AVDD.n927 AVDD.n926 185
R5994 AVDD.n929 AVDD.n796 185
R5995 AVDD.n932 AVDD.n931 185
R5996 AVDD.n793 AVDD.n792 185
R5997 AVDD.n938 AVDD.n937 185
R5998 AVDD.n941 AVDD.n940 185
R5999 AVDD.n791 AVDD.n786 185
R6000 AVDD.n949 AVDD.n948 185
R6001 AVDD.n966 AVDD.n965 185
R6002 AVDD.n963 AVDD.n783 185
R6003 AVDD.n962 AVDD.n950 185
R6004 AVDD.n960 AVDD.n959 185
R6005 AVDD.n955 AVDD.n952 185
R6006 AVDD.n779 AVDD.n778 185
R6007 AVDD.n976 AVDD.n975 185
R6008 AVDD.n977 AVDD.n976 185
R6009 AVDD.n780 AVDD.n769 185
R6010 AVDD.n777 AVDD.n769 185
R6011 AVDD.n988 AVDD.n987 185
R6012 AVDD.n987 AVDD.n986 185
R6013 AVDD.n989 AVDD.n764 185
R6014 AVDD.n764 AVDD.n763 185
R6015 AVDD.n998 AVDD.n997 185
R6016 AVDD.n999 AVDD.n998 185
R6017 AVDD.n766 AVDD.n755 185
R6018 AVDD.n756 AVDD.n755 185
R6019 AVDD.n1023 AVDD.n1022 185
R6020 AVDD.n1022 AVDD.n1021 185
R6021 AVDD.n752 AVDD.n751 185
R6022 AVDD.n1020 AVDD.n751 185
R6023 AVDD.n1033 AVDD.n1032 185
R6024 AVDD.n1034 AVDD.n1033 185
R6025 AVDD.n739 AVDD.n737 185
R6026 AVDD.n741 AVDD.n739 185
R6027 AVDD.n1064 AVDD.n1063 185
R6028 AVDD.n1063 AVDD.n1062 185
R6029 AVDD.n1051 AVDD.n740 185
R6030 AVDD.n1061 AVDD.n740 185
R6031 AVDD.n1059 AVDD.n1058 185
R6032 AVDD.n1060 AVDD.n1059 185
R6033 AVDD.n1057 AVDD.n731 185
R6034 AVDD.n731 AVDD.n730 185
R6035 AVDD.n1077 AVDD.n1076 185
R6036 AVDD.n1078 AVDD.n1077 185
R6037 AVDD.n733 AVDD.n719 185
R6038 AVDD.n1079 AVDD.n719 185
R6039 AVDD.n1096 AVDD.n1095 185
R6040 AVDD.n1095 AVDD.n1094 185
R6041 AVDD.n720 AVDD.n716 185
R6042 AVDD.n1093 AVDD.n720 185
R6043 AVDD.n1101 AVDD.n706 185
R6044 AVDD.n708 AVDD.n706 185
R6045 AVDD.n1112 AVDD.n707 185
R6046 AVDD.n1112 AVDD.n1111 185
R6047 AVDD.n1114 AVDD.n1113 185
R6048 AVDD.n1113 AVDD.n689 185
R6049 AVDD.n1116 AVDD.n687 185
R6050 AVDD.n1122 AVDD.n687 185
R6051 AVDD.n1124 AVDD.n688 185
R6052 AVDD.n1124 AVDD.n1123 185
R6053 AVDD.n1125 AVDD.n683 185
R6054 AVDD.n1126 AVDD.n1125 185
R6055 AVDD.n1133 AVDD.n682 185
R6056 AVDD.n682 AVDD.n594 185
R6057 AVDD.n1135 AVDD.n1134 185
R6058 AVDD.n681 AVDD.n680 185
R6059 AVDD.n679 AVDD.n678 185
R6060 AVDD.n1137 AVDD.n679 185
R6061 AVDD.n677 AVDD.n676 185
R6062 AVDD.n597 AVDD.n596 185
R6063 AVDD.n599 AVDD.n598 185
R6064 AVDD.n602 AVDD.n601 185
R6065 AVDD.n604 AVDD.n603 185
R6066 AVDD.n607 AVDD.n606 185
R6067 AVDD.n609 AVDD.n608 185
R6068 AVDD.n613 AVDD.n612 185
R6069 AVDD.n615 AVDD.n614 185
R6070 AVDD.n617 AVDD.n616 185
R6071 AVDD.n619 AVDD.n618 185
R6072 AVDD.n622 AVDD.n621 185
R6073 AVDD.n624 AVDD.n623 185
R6074 AVDD.n627 AVDD.n626 185
R6075 AVDD.n629 AVDD.n628 185
R6076 AVDD.n632 AVDD.n631 185
R6077 AVDD.n634 AVDD.n633 185
R6078 AVDD.n637 AVDD.n636 185
R6079 AVDD.n639 AVDD.n638 185
R6080 AVDD.n642 AVDD.n641 185
R6081 AVDD.n644 AVDD.n643 185
R6082 AVDD.n647 AVDD.n646 185
R6083 AVDD.n649 AVDD.n648 185
R6084 AVDD.n652 AVDD.n651 185
R6085 AVDD.n654 AVDD.n653 185
R6086 AVDD.n658 AVDD.n657 185
R6087 AVDD.n660 AVDD.n659 185
R6088 AVDD.n662 AVDD.n661 185
R6089 AVDD.n664 AVDD.n663 185
R6090 AVDD.n667 AVDD.n666 185
R6091 AVDD.n669 AVDD.n668 185
R6092 AVDD.n672 AVDD.n671 185
R6093 AVDD.n674 AVDD.n673 185
R6094 AVDD.n592 AVDD.n590 185
R6095 AVDD.n1139 AVDD.n1138 185
R6096 AVDD.n1138 AVDD.n1137 185
R6097 AVDD.n593 AVDD.n591 185
R6098 AVDD.n594 AVDD.n593 185
R6099 AVDD.n1128 AVDD.n1127 185
R6100 AVDD.n1127 AVDD.n1126 185
R6101 AVDD.n692 AVDD.n686 185
R6102 AVDD.n1123 AVDD.n686 185
R6103 AVDD.n1121 AVDD.n1120 185
R6104 AVDD.n1122 AVDD.n1121 185
R6105 AVDD.n711 AVDD.n690 185
R6106 AVDD.n690 AVDD.n689 185
R6107 AVDD.n1110 AVDD.n1109 185
R6108 AVDD.n1111 AVDD.n1110 185
R6109 AVDD.n723 AVDD.n709 185
R6110 AVDD.n709 AVDD.n708 185
R6111 AVDD.n1092 AVDD.n1091 185
R6112 AVDD.n1093 AVDD.n1092 185
R6113 AVDD.n727 AVDD.n721 185
R6114 AVDD.n1094 AVDD.n721 185
R6115 AVDD.n1081 AVDD.n1080 185
R6116 AVDD.n1080 AVDD.n1079 185
R6117 AVDD.n729 AVDD.n726 185
R6118 AVDD.n1078 AVDD.n729 185
R6119 AVDD.n1048 AVDD.n744 185
R6120 AVDD.n744 AVDD.n730 185
R6121 AVDD.n1050 AVDD.n1049 185
R6122 AVDD.n1060 AVDD.n1050 185
R6123 AVDD.n1040 AVDD.n743 185
R6124 AVDD.n1061 AVDD.n743 185
R6125 AVDD.n1039 AVDD.n742 185
R6126 AVDD.n1062 AVDD.n742 185
R6127 AVDD.n1037 AVDD.n1036 185
R6128 AVDD.n1036 AVDD.n741 185
R6129 AVDD.n1035 AVDD.n750 185
R6130 AVDD.n1035 AVDD.n1034 185
R6131 AVDD.n759 AVDD.n749 185
R6132 AVDD.n1020 AVDD.n749 185
R6133 AVDD.n1019 AVDD.n1018 185
R6134 AVDD.n1021 AVDD.n1019 185
R6135 AVDD.n1002 AVDD.n757 185
R6136 AVDD.n757 AVDD.n756 185
R6137 AVDD.n1001 AVDD.n1000 185
R6138 AVDD.n1000 AVDD.n999 185
R6139 AVDD.n772 AVDD.n762 185
R6140 AVDD.n763 AVDD.n762 185
R6141 AVDD.n985 AVDD.n984 185
R6142 AVDD.n986 AVDD.n985 185
R6143 AVDD.n980 AVDD.n770 185
R6144 AVDD.n777 AVDD.n770 185
R6145 AVDD.n979 AVDD.n978 185
R6146 AVDD.n978 AVDD.n977 185
R6147 AVDD.n1746 AVDD.n1745 128.922
R6148 AVDD.n1747 AVDD.n1746 128.922
R6149 AVDD.n495 AVDD.n490 115.954
R6150 AVDD.n518 AVDD.t323 113.576
R6151 AVDD.n527 AVDD.t185 113.576
R6152 AVDD.n1165 AVDD.t360 113.576
R6153 AVDD.n1174 AVDD.t133 113.576
R6154 AVDD.n1763 AVDD.t306 113.576
R6155 AVDD.n1752 AVDD.t155 113.576
R6156 AVDD.n211 AVDD.t174 113.576
R6157 AVDD.n225 AVDD.t336 113.576
R6158 AVDD.n250 AVDD.t158 113.576
R6159 AVDD.n259 AVDD.t320 113.576
R6160 AVDD.n290 AVDD.t213 113.576
R6161 AVDD.n301 AVDD.t331 113.576
R6162 AVDD.n352 AVDD.t161 113.576
R6163 AVDD.n2934 AVDD.t314 113.576
R6164 AVDD.n420 AVDD.t243 113.576
R6165 AVDD.n429 AVDD.t366 113.576
R6166 AVDD.n483 AVDD.t352 113.576
R6167 AVDD.n794 AVDD.t201 113.576
R6168 AVDD.n795 AVDD.t300 113.576
R6169 AVDD.n903 AVDD.t346 113.576
R6170 AVDD.n820 AVDD.t129 113.576
R6171 AVDD.n841 AVDD.t260 113.576
R6172 AVDD.n842 AVDD.t393 113.576
R6173 AVDD.n105 AVDD.t226 113.576
R6174 AVDD.n3270 AVDD.t407 113.576
R6175 AVDD.n142 AVDD.t265 113.576
R6176 AVDD.n147 AVDD.t339 113.576
R6177 AVDD.n173 AVDD.t204 113.576
R6178 AVDD.n178 AVDD.t363 113.576
R6179 AVDD.n1356 AVDD.t398 113.576
R6180 AVDD.n1369 AVDD.t240 113.576
R6181 AVDD.n1396 AVDD.t372 113.576
R6182 AVDD.n1663 AVDD.t218 113.576
R6183 AVDD.n1442 AVDD.t191 113.576
R6184 AVDD.n1445 AVDD.t311 113.576
R6185 AVDD.n1497 AVDD.t375 113.576
R6186 AVDD.n1545 AVDD.t317 113.576
R6187 AVDD.n2260 AVDD.t246 113.576
R6188 AVDD.n2226 AVDD.t369 113.576
R6189 AVDD.n2188 AVDD.t355 113.576
R6190 AVDD.n518 AVDD.t334 113.576
R6191 AVDD.n527 AVDD.t199 113.576
R6192 AVDD.n1165 AVDD.t378 113.576
R6193 AVDD.n1174 AVDD.t146 113.576
R6194 AVDD.n1763 AVDD.t309 113.576
R6195 AVDD.n1752 AVDD.t164 113.576
R6196 AVDD.n211 AVDD.t180 113.576
R6197 AVDD.n225 AVDD.t342 113.576
R6198 AVDD.n250 AVDD.t168 113.576
R6199 AVDD.n259 AVDD.t329 113.576
R6200 AVDD.n290 AVDD.t283 113.576
R6201 AVDD.n301 AVDD.t417 113.576
R6202 AVDD.n352 AVDD.t170 113.576
R6203 AVDD.n2934 AVDD.t231 113.576
R6204 AVDD.n420 AVDD.t140 113.576
R6205 AVDD.n429 AVDD.t281 113.576
R6206 AVDD.n483 AVDD.t268 113.576
R6207 AVDD.n105 AVDD.t235 113.576
R6208 AVDD.n3270 AVDD.t415 113.576
R6209 AVDD.n142 AVDD.t276 113.576
R6210 AVDD.n147 AVDD.t344 113.576
R6211 AVDD.n173 AVDD.t209 113.576
R6212 AVDD.n178 AVDD.t380 113.576
R6213 AVDD.n1356 AVDD.t403 113.576
R6214 AVDD.n1369 AVDD.t251 113.576
R6215 AVDD.n1396 AVDD.t386 113.576
R6216 AVDD.n1663 AVDD.t229 113.576
R6217 AVDD.n1442 AVDD.t270 113.576
R6218 AVDD.n1445 AVDD.t401 113.576
R6219 AVDD.n1497 AVDD.t391 113.576
R6220 AVDD.n1545 AVDD.t233 113.576
R6221 AVDD.n2260 AVDD.t143 113.576
R6222 AVDD.n2226 AVDD.t285 113.576
R6223 AVDD.n2188 AVDD.t274 113.576
R6224 AVDD.n1894 AVDD.n511 105.788
R6225 AVDD.n2617 AVDD.t388 102.6
R6226 AVDD.n2344 AVDD.t287 102.6
R6227 AVDD.n2589 AVDD.t195 102.6
R6228 AVDD.n2572 AVDD.t253 102.6
R6229 AVDD.n2551 AVDD.t188 102.6
R6230 AVDD.n2529 AVDD.t207 102.6
R6231 AVDD.n2482 AVDD.t396 102.6
R6232 AVDD.n2495 AVDD.t405 102.6
R6233 AVDD.n2505 AVDD.t298 102.6
R6234 AVDD.n2513 AVDD.t216 102.6
R6235 AVDD.n2436 AVDD.t293 102.6
R6236 AVDD.n2379 AVDD.t211 102.6
R6237 AVDD.n2413 AVDD.t221 102.6
R6238 AVDD.n2395 AVDD.t410 102.6
R6239 AVDD.n703 AVDD.t303 102.6
R6240 AVDD.n694 AVDD.t349 102.6
R6241 AVDD.n701 AVDD.t148 102.6
R6242 AVDD.n695 AVDD.t182 102.6
R6243 AVDD.n700 AVDD.t278 102.6
R6244 AVDD.n696 AVDD.t412 102.6
R6245 AVDD.n699 AVDD.t223 102.6
R6246 AVDD.n1072 AVDD.t326 102.6
R6247 AVDD.n1053 AVDD.t263 102.6
R6248 AVDD.n1027 AVDD.t272 102.6
R6249 AVDD.n970 AVDD.t152 102.6
R6250 AVDD.n1085 AVDD.t257 102.6
R6251 AVDD.n1044 AVDD.t166 102.6
R6252 AVDD.n1014 AVDD.t172 102.6
R6253 AVDD.n2154 AVDD.t237 102.6
R6254 AVDD.n2136 AVDD.t249 102.6
R6255 AVDD.n2684 AVDD.t255 102.6
R6256 AVDD.n2698 AVDD.t382 102.6
R6257 AVDD.n2085 AVDD.t137 102.6
R6258 AVDD.n2063 AVDD.t384 102.6
R6259 AVDD.n2735 AVDD.t358 102.6
R6260 AVDD.n2748 AVDD.t289 102.6
R6261 AVDD.n2762 AVDD.t291 102.6
R6262 AVDD.n2015 AVDD.t296 102.6
R6263 AVDD.n2787 AVDD.t177 102.6
R6264 AVDD.n2799 AVDD.t197 102.6
R6265 AVDD.n2813 AVDD.t127 102.6
R6266 AVDD.n1951 AVDD.t419 102.6
R6267 AVDD.n979 AVDD.n774 101.272
R6268 AVDD.n2321 AVDD.n2187 100.141
R6269 AVDD.n975 AVDD.n779 95.624
R6270 AVDD.n294 AVDD.n62 95.2946
R6271 AVDD.n2999 AVDD.n295 95.2946
R6272 AVDD.n1139 AVDD.n591 90.3534
R6273 AVDD.n2175 AVDD.n98 89.977
R6274 AVDD.n1134 AVDD.n1133 84.7064
R6275 AVDD.n1735 AVDD.n1734 81.177
R6276 AVDD.n1733 AVDD.n42 81.177
R6277 AVDD.n2992 AVDD.n304 72.7879
R6278 AVDD.n2990 AVDD.n2989 72.7879
R6279 AVDD.n318 AVDD.n317 72.7879
R6280 AVDD.n2978 AVDD.n2977 72.7879
R6281 AVDD.n2970 AVDD.n323 72.7879
R6282 AVDD.n2968 AVDD.n2967 72.7879
R6283 AVDD.n2960 AVDD.n332 72.7879
R6284 AVDD.n2958 AVDD.n2957 72.7879
R6285 AVDD.n2950 AVDD.n340 72.7879
R6286 AVDD.n2948 AVDD.n2947 72.7879
R6287 AVDD.n357 AVDD.n356 72.7879
R6288 AVDD.n2939 AVDD.n2938 72.7879
R6289 AVDD.n2930 AVDD.n362 72.7879
R6290 AVDD.n2928 AVDD.n2927 72.7879
R6291 AVDD.n2920 AVDD.n376 72.7879
R6292 AVDD.n2918 AVDD.n2917 72.7879
R6293 AVDD.n2910 AVDD.n398 72.7879
R6294 AVDD.n2908 AVDD.n2907 72.7879
R6295 AVDD.n2900 AVDD.n407 72.7879
R6296 AVDD.n2898 AVDD.n2897 72.7879
R6297 AVDD.n2886 AVDD.n415 72.7879
R6298 AVDD.n2884 AVDD.n2883 72.7879
R6299 AVDD.n2876 AVDD.n424 72.7879
R6300 AVDD.n2874 AVDD.n2873 72.7879
R6301 AVDD.n440 AVDD.n439 72.7879
R6302 AVDD.n2862 AVDD.n2861 72.7879
R6303 AVDD.n2854 AVDD.n445 72.7879
R6304 AVDD.n2852 AVDD.n2851 72.7879
R6305 AVDD.n455 AVDD.n454 72.7879
R6306 AVDD.n2843 AVDD.n2842 72.7879
R6307 AVDD.n497 AVDD.n491 72.7879
R6308 AVDD.n1333 AVDD.n43 72.7879
R6309 AVDD.n1348 AVDD.n44 72.7879
R6310 AVDD.n1351 AVDD.n45 72.7879
R6311 AVDD.n1361 AVDD.n46 72.7879
R6312 AVDD.n1364 AVDD.n47 72.7879
R6313 AVDD.n1374 AVDD.n48 72.7879
R6314 AVDD.n1377 AVDD.n49 72.7879
R6315 AVDD.n1389 AVDD.n50 72.7879
R6316 AVDD.n1697 AVDD.n51 72.7879
R6317 AVDD.n1690 AVDD.n52 72.7879
R6318 AVDD.n1679 AVDD.n53 72.7879
R6319 AVDD.n1672 AVDD.n54 72.7879
R6320 AVDD.n1667 AVDD.n55 72.7879
R6321 AVDD.n1659 AVDD.n56 72.7879
R6322 AVDD.n1654 AVDD.n57 72.7879
R6323 AVDD.n1647 AVDD.n58 72.7879
R6324 AVDD.n1640 AVDD.n59 72.7879
R6325 AVDD.n1635 AVDD.n60 72.7879
R6326 AVDD.n1624 AVDD.n61 72.7879
R6327 AVDD.n1613 AVDD.n63 72.7879
R6328 AVDD.n1450 AVDD.n64 72.7879
R6329 AVDD.n1606 AVDD.n65 72.7879
R6330 AVDD.n1599 AVDD.n66 72.7879
R6331 AVDD.n1594 AVDD.n67 72.7879
R6332 AVDD.n1587 AVDD.n68 72.7879
R6333 AVDD.n1580 AVDD.n69 72.7879
R6334 AVDD.n1575 AVDD.n70 72.7879
R6335 AVDD.n1568 AVDD.n71 72.7879
R6336 AVDD.n1557 AVDD.n72 72.7879
R6337 AVDD.n1501 AVDD.n73 72.7879
R6338 AVDD.n1549 AVDD.n74 72.7879
R6339 AVDD.n1541 AVDD.n75 72.7879
R6340 AVDD.n1536 AVDD.n76 72.7879
R6341 AVDD.n1529 AVDD.n77 72.7879
R6342 AVDD.n1524 AVDD.n78 72.7879
R6343 AVDD.n3298 AVDD.n12 72.7879
R6344 AVDD.n79 AVDD.n11 72.7879
R6345 AVDD.n2240 AVDD.n80 72.7879
R6346 AVDD.n2242 AVDD.n81 72.7879
R6347 AVDD.n2254 AVDD.n82 72.7879
R6348 AVDD.n2265 AVDD.n83 72.7879
R6349 AVDD.n2268 AVDD.n84 72.7879
R6350 AVDD.n2275 AVDD.n85 72.7879
R6351 AVDD.n2291 AVDD.n86 72.7879
R6352 AVDD.n2294 AVDD.n87 72.7879
R6353 AVDD.n2304 AVDD.n88 72.7879
R6354 AVDD.n2307 AVDD.n89 72.7879
R6355 AVDD.n2316 AVDD.n90 72.7879
R6356 AVDD.n2328 AVDD.n91 72.7879
R6357 AVDD.n1891 AVDD.n1890 72.7879
R6358 AVDD.n1879 AVDD.n520 72.7879
R6359 AVDD.n1877 AVDD.n1876 72.7879
R6360 AVDD.n531 AVDD.n530 72.7879
R6361 AVDD.n1868 AVDD.n1867 72.7879
R6362 AVDD.n544 AVDD.n543 72.7879
R6363 AVDD.n1856 AVDD.n1855 72.7879
R6364 AVDD.n1848 AVDD.n549 72.7879
R6365 AVDD.n1846 AVDD.n1845 72.7879
R6366 AVDD.n1837 AVDD.n1144 72.7879
R6367 AVDD.n1835 AVDD.n1834 72.7879
R6368 AVDD.n1159 AVDD.n1158 72.7879
R6369 AVDD.n1823 AVDD.n1822 72.7879
R6370 AVDD.n1820 AVDD.n1819 72.7879
R6371 AVDD.n1812 AVDD.n1169 72.7879
R6372 AVDD.n1810 AVDD.n1809 72.7879
R6373 AVDD.n1185 AVDD.n1184 72.7879
R6374 AVDD.n1798 AVDD.n1797 72.7879
R6375 AVDD.n1790 AVDD.n1190 72.7879
R6376 AVDD.n1788 AVDD.n1787 72.7879
R6377 AVDD.n1780 AVDD.n1199 72.7879
R6378 AVDD.n1778 AVDD.n1777 72.7879
R6379 AVDD.n1770 AVDD.n1205 72.7879
R6380 AVDD.n1768 AVDD.n1767 72.7879
R6381 AVDD.n1759 AVDD.n1219 72.7879
R6382 AVDD.n1757 AVDD.n1756 72.7879
R6383 AVDD.n1748 AVDD.n1227 72.7879
R6384 AVDD.n1738 AVDD.n1729 72.7879
R6385 AVDD.n1736 AVDD.n1735 72.7879
R6386 AVDD.n3103 AVDD.n198 72.7879
R6387 AVDD.n3101 AVDD.n3100 72.7879
R6388 AVDD.n3093 AVDD.n213 72.7879
R6389 AVDD.n3091 AVDD.n3090 72.7879
R6390 AVDD.n3083 AVDD.n220 72.7879
R6391 AVDD.n3081 AVDD.n3080 72.7879
R6392 AVDD.n236 AVDD.n235 72.7879
R6393 AVDD.n3069 AVDD.n3068 72.7879
R6394 AVDD.n3061 AVDD.n242 72.7879
R6395 AVDD.n3059 AVDD.n3058 72.7879
R6396 AVDD.n3047 AVDD.n252 72.7879
R6397 AVDD.n3045 AVDD.n3044 72.7879
R6398 AVDD.n263 AVDD.n262 72.7879
R6399 AVDD.n3036 AVDD.n3035 72.7879
R6400 AVDD.n276 AVDD.n275 72.7879
R6401 AVDD.n3024 AVDD.n3023 72.7879
R6402 AVDD.n3016 AVDD.n282 72.7879
R6403 AVDD.n3014 AVDD.n3013 72.7879
R6404 AVDD.n3002 AVDD.n292 72.7879
R6405 AVDD.n3000 AVDD.n2999 72.7879
R6406 AVDD.n3296 AVDD.n3295 72.7879
R6407 AVDD.n3285 AVDD.n14 72.7879
R6408 AVDD.n3279 AVDD.n15 72.7879
R6409 AVDD.n3274 AVDD.n16 72.7879
R6410 AVDD.n3266 AVDD.n17 72.7879
R6411 AVDD.n3261 AVDD.n18 72.7879
R6412 AVDD.n3254 AVDD.n19 72.7879
R6413 AVDD.n3249 AVDD.n20 72.7879
R6414 AVDD.n3242 AVDD.n21 72.7879
R6415 AVDD.n3235 AVDD.n22 72.7879
R6416 AVDD.n3230 AVDD.n23 72.7879
R6417 AVDD.n138 AVDD.n24 72.7879
R6418 AVDD.n3219 AVDD.n25 72.7879
R6419 AVDD.n3214 AVDD.n26 72.7879
R6420 AVDD.n3207 AVDD.n27 72.7879
R6421 AVDD.n3202 AVDD.n28 72.7879
R6422 AVDD.n156 AVDD.n29 72.7879
R6423 AVDD.n3191 AVDD.n30 72.7879
R6424 AVDD.n3184 AVDD.n31 72.7879
R6425 AVDD.n3179 AVDD.n32 72.7879
R6426 AVDD.n3172 AVDD.n33 72.7879
R6427 AVDD.n3167 AVDD.n34 72.7879
R6428 AVDD.n3160 AVDD.n35 72.7879
R6429 AVDD.n3149 AVDD.n36 72.7879
R6430 AVDD.n3144 AVDD.n37 72.7879
R6431 AVDD.n3137 AVDD.n38 72.7879
R6432 AVDD.n3132 AVDD.n39 72.7879
R6433 AVDD.n3122 AVDD.n40 72.7879
R6434 AVDD.n3117 AVDD.n41 72.7879
R6435 AVDD.n3296 AVDD.n96 72.7879
R6436 AVDD.n3278 AVDD.n14 72.7879
R6437 AVDD.n3275 AVDD.n15 72.7879
R6438 AVDD.n3265 AVDD.n16 72.7879
R6439 AVDD.n3262 AVDD.n17 72.7879
R6440 AVDD.n3253 AVDD.n18 72.7879
R6441 AVDD.n3250 AVDD.n19 72.7879
R6442 AVDD.n3241 AVDD.n20 72.7879
R6443 AVDD.n3234 AVDD.n21 72.7879
R6444 AVDD.n3231 AVDD.n22 72.7879
R6445 AVDD.n137 AVDD.n23 72.7879
R6446 AVDD.n3220 AVDD.n24 72.7879
R6447 AVDD.n3215 AVDD.n25 72.7879
R6448 AVDD.n3206 AVDD.n26 72.7879
R6449 AVDD.n3203 AVDD.n27 72.7879
R6450 AVDD.n155 AVDD.n28 72.7879
R6451 AVDD.n3192 AVDD.n29 72.7879
R6452 AVDD.n3183 AVDD.n30 72.7879
R6453 AVDD.n3180 AVDD.n31 72.7879
R6454 AVDD.n3171 AVDD.n32 72.7879
R6455 AVDD.n3168 AVDD.n33 72.7879
R6456 AVDD.n3159 AVDD.n34 72.7879
R6457 AVDD.n3148 AVDD.n35 72.7879
R6458 AVDD.n3145 AVDD.n36 72.7879
R6459 AVDD.n3136 AVDD.n37 72.7879
R6460 AVDD.n3133 AVDD.n38 72.7879
R6461 AVDD.n3121 AVDD.n39 72.7879
R6462 AVDD.n3118 AVDD.n40 72.7879
R6463 AVDD.n187 AVDD.n41 72.7879
R6464 AVDD.n1347 AVDD.n43 72.7879
R6465 AVDD.n1352 AVDD.n44 72.7879
R6466 AVDD.n1360 AVDD.n45 72.7879
R6467 AVDD.n1365 AVDD.n46 72.7879
R6468 AVDD.n1373 AVDD.n47 72.7879
R6469 AVDD.n1378 AVDD.n48 72.7879
R6470 AVDD.n1388 AVDD.n49 72.7879
R6471 AVDD.n1698 AVDD.n50 72.7879
R6472 AVDD.n1689 AVDD.n51 72.7879
R6473 AVDD.n1678 AVDD.n52 72.7879
R6474 AVDD.n1671 AVDD.n53 72.7879
R6475 AVDD.n1668 AVDD.n54 72.7879
R6476 AVDD.n1658 AVDD.n55 72.7879
R6477 AVDD.n1655 AVDD.n56 72.7879
R6478 AVDD.n1646 AVDD.n57 72.7879
R6479 AVDD.n1639 AVDD.n58 72.7879
R6480 AVDD.n1636 AVDD.n59 72.7879
R6481 AVDD.n1623 AVDD.n60 72.7879
R6482 AVDD.n1443 AVDD.n61 72.7879
R6483 AVDD.n1449 AVDD.n63 72.7879
R6484 AVDD.n1607 AVDD.n64 72.7879
R6485 AVDD.n1598 AVDD.n65 72.7879
R6486 AVDD.n1595 AVDD.n66 72.7879
R6487 AVDD.n1586 AVDD.n67 72.7879
R6488 AVDD.n1579 AVDD.n68 72.7879
R6489 AVDD.n1576 AVDD.n69 72.7879
R6490 AVDD.n1567 AVDD.n70 72.7879
R6491 AVDD.n1556 AVDD.n71 72.7879
R6492 AVDD.n1500 AVDD.n72 72.7879
R6493 AVDD.n1550 AVDD.n73 72.7879
R6494 AVDD.n1540 AVDD.n74 72.7879
R6495 AVDD.n1537 AVDD.n75 72.7879
R6496 AVDD.n1528 AVDD.n76 72.7879
R6497 AVDD.n1525 AVDD.n77 72.7879
R6498 AVDD.n1518 AVDD.n78 72.7879
R6499 AVDD.n3299 AVDD.n3298 72.7879
R6500 AVDD.n2239 AVDD.n79 72.7879
R6501 AVDD.n2243 AVDD.n80 72.7879
R6502 AVDD.n2255 AVDD.n81 72.7879
R6503 AVDD.n2264 AVDD.n82 72.7879
R6504 AVDD.n2269 AVDD.n83 72.7879
R6505 AVDD.n2276 AVDD.n84 72.7879
R6506 AVDD.n2290 AVDD.n85 72.7879
R6507 AVDD.n2295 AVDD.n86 72.7879
R6508 AVDD.n2303 AVDD.n87 72.7879
R6509 AVDD.n2308 AVDD.n88 72.7879
R6510 AVDD.n2315 AVDD.n89 72.7879
R6511 AVDD.n2327 AVDD.n90 72.7879
R6512 AVDD.n2324 AVDD.n91 72.7879
R6513 AVDD.n491 AVDD.n456 72.7879
R6514 AVDD.n2844 AVDD.n2843 72.7879
R6515 AVDD.n454 AVDD.n447 72.7879
R6516 AVDD.n2853 AVDD.n2852 72.7879
R6517 AVDD.n445 AVDD.n441 72.7879
R6518 AVDD.n2863 AVDD.n2862 72.7879
R6519 AVDD.n439 AVDD.n426 72.7879
R6520 AVDD.n2875 AVDD.n2874 72.7879
R6521 AVDD.n424 AVDD.n417 72.7879
R6522 AVDD.n2885 AVDD.n2884 72.7879
R6523 AVDD.n415 AVDD.n409 72.7879
R6524 AVDD.n2899 AVDD.n2898 72.7879
R6525 AVDD.n407 AVDD.n400 72.7879
R6526 AVDD.n2909 AVDD.n2908 72.7879
R6527 AVDD.n398 AVDD.n378 72.7879
R6528 AVDD.n2919 AVDD.n2918 72.7879
R6529 AVDD.n376 AVDD.n364 72.7879
R6530 AVDD.n2929 AVDD.n2928 72.7879
R6531 AVDD.n362 AVDD.n358 72.7879
R6532 AVDD.n2940 AVDD.n2939 72.7879
R6533 AVDD.n356 AVDD.n342 72.7879
R6534 AVDD.n2949 AVDD.n2948 72.7879
R6535 AVDD.n340 AVDD.n334 72.7879
R6536 AVDD.n2959 AVDD.n2958 72.7879
R6537 AVDD.n332 AVDD.n325 72.7879
R6538 AVDD.n2969 AVDD.n2968 72.7879
R6539 AVDD.n323 AVDD.n319 72.7879
R6540 AVDD.n2979 AVDD.n2978 72.7879
R6541 AVDD.n317 AVDD.n306 72.7879
R6542 AVDD.n2991 AVDD.n2990 72.7879
R6543 AVDD.n304 AVDD.n303 72.7879
R6544 AVDD.n3001 AVDD.n3000 72.7879
R6545 AVDD.n292 AVDD.n284 72.7879
R6546 AVDD.n3015 AVDD.n3014 72.7879
R6547 AVDD.n282 AVDD.n277 72.7879
R6548 AVDD.n3025 AVDD.n3024 72.7879
R6549 AVDD.n275 AVDD.n264 72.7879
R6550 AVDD.n3037 AVDD.n3036 72.7879
R6551 AVDD.n262 AVDD.n254 72.7879
R6552 AVDD.n3046 AVDD.n3045 72.7879
R6553 AVDD.n252 AVDD.n244 72.7879
R6554 AVDD.n3060 AVDD.n3059 72.7879
R6555 AVDD.n242 AVDD.n237 72.7879
R6556 AVDD.n3070 AVDD.n3069 72.7879
R6557 AVDD.n235 AVDD.n222 72.7879
R6558 AVDD.n3082 AVDD.n3081 72.7879
R6559 AVDD.n220 AVDD.n215 72.7879
R6560 AVDD.n3092 AVDD.n3091 72.7879
R6561 AVDD.n213 AVDD.n201 72.7879
R6562 AVDD.n3102 AVDD.n3101 72.7879
R6563 AVDD.n1732 AVDD.n198 72.7879
R6564 AVDD.n1737 AVDD.n1736 72.7879
R6565 AVDD.n1729 AVDD.n1229 72.7879
R6566 AVDD.n1227 AVDD.n1221 72.7879
R6567 AVDD.n1758 AVDD.n1757 72.7879
R6568 AVDD.n1219 AVDD.n1207 72.7879
R6569 AVDD.n1769 AVDD.n1768 72.7879
R6570 AVDD.n1205 AVDD.n1201 72.7879
R6571 AVDD.n1779 AVDD.n1778 72.7879
R6572 AVDD.n1199 AVDD.n1192 72.7879
R6573 AVDD.n1789 AVDD.n1788 72.7879
R6574 AVDD.n1190 AVDD.n1186 72.7879
R6575 AVDD.n1799 AVDD.n1798 72.7879
R6576 AVDD.n1184 AVDD.n1171 72.7879
R6577 AVDD.n1811 AVDD.n1810 72.7879
R6578 AVDD.n1169 AVDD.n1162 72.7879
R6579 AVDD.n1821 AVDD.n1820 72.7879
R6580 AVDD.n1824 AVDD.n1823 72.7879
R6581 AVDD.n1158 AVDD.n1146 72.7879
R6582 AVDD.n1836 AVDD.n1835 72.7879
R6583 AVDD.n1144 AVDD.n551 72.7879
R6584 AVDD.n1847 AVDD.n1846 72.7879
R6585 AVDD.n549 AVDD.n545 72.7879
R6586 AVDD.n1857 AVDD.n1856 72.7879
R6587 AVDD.n543 AVDD.n532 72.7879
R6588 AVDD.n1869 AVDD.n1868 72.7879
R6589 AVDD.n530 AVDD.n522 72.7879
R6590 AVDD.n1878 AVDD.n1877 72.7879
R6591 AVDD.n520 AVDD.n513 72.7879
R6592 AVDD.n1892 AVDD.n1891 72.7879
R6593 AVDD.n1136 AVDD.n1135 72.7879
R6594 AVDD.n677 AVDD.n595 72.7879
R6595 AVDD.n600 AVDD.n599 72.7879
R6596 AVDD.n605 AVDD.n604 72.7879
R6597 AVDD.n610 AVDD.n609 72.7879
R6598 AVDD.n614 AVDD.n611 72.7879
R6599 AVDD.n620 AVDD.n619 72.7879
R6600 AVDD.n625 AVDD.n624 72.7879
R6601 AVDD.n630 AVDD.n629 72.7879
R6602 AVDD.n635 AVDD.n634 72.7879
R6603 AVDD.n640 AVDD.n639 72.7879
R6604 AVDD.n645 AVDD.n644 72.7879
R6605 AVDD.n650 AVDD.n649 72.7879
R6606 AVDD.n655 AVDD.n654 72.7879
R6607 AVDD.n659 AVDD.n656 72.7879
R6608 AVDD.n665 AVDD.n664 72.7879
R6609 AVDD.n670 AVDD.n669 72.7879
R6610 AVDD.n675 AVDD.n674 72.7879
R6611 AVDD.n951 AVDD.n778 72.7879
R6612 AVDD.n961 AVDD.n960 72.7879
R6613 AVDD.n964 AVDD.n963 72.7879
R6614 AVDD.n949 AVDD.n785 72.7879
R6615 AVDD.n940 AVDD.n939 72.7879
R6616 AVDD.n930 AVDD.n792 72.7879
R6617 AVDD.n929 AVDD.n928 72.7879
R6618 AVDD.n917 AVDD.n797 72.7879
R6619 AVDD.n916 AVDD.n805 72.7879
R6620 AVDD.n909 AVDD.n908 72.7879
R6621 AVDD.n898 AVDD.n810 72.7879
R6622 AVDD.n897 AVDD.n818 72.7879
R6623 AVDD.n890 AVDD.n889 72.7879
R6624 AVDD.n880 AVDD.n824 72.7879
R6625 AVDD.n879 AVDD.n832 72.7879
R6626 AVDD.n869 AVDD.n868 72.7879
R6627 AVDD.n866 AVDD.n839 72.7879
R6628 AVDD.n859 AVDD.n858 72.7879
R6629 AVDD.n846 AVDD.n845 72.7879
R6630 AVDD.n845 AVDD.n775 72.7879
R6631 AVDD.n858 AVDD.n857 72.7879
R6632 AVDD.n844 AVDD.n839 72.7879
R6633 AVDD.n870 AVDD.n869 72.7879
R6634 AVDD.n867 AVDD.n832 72.7879
R6635 AVDD.n881 AVDD.n880 72.7879
R6636 AVDD.n889 AVDD.n888 72.7879
R6637 AVDD.n823 AVDD.n818 72.7879
R6638 AVDD.n899 AVDD.n898 72.7879
R6639 AVDD.n908 AVDD.n907 72.7879
R6640 AVDD.n809 AVDD.n805 72.7879
R6641 AVDD.n918 AVDD.n917 72.7879
R6642 AVDD.n928 AVDD.n927 72.7879
R6643 AVDD.n931 AVDD.n930 72.7879
R6644 AVDD.n939 AVDD.n938 72.7879
R6645 AVDD.n791 AVDD.n785 72.7879
R6646 AVDD.n965 AVDD.n964 72.7879
R6647 AVDD.n962 AVDD.n961 72.7879
R6648 AVDD.n952 AVDD.n951 72.7879
R6649 AVDD.n1136 AVDD.n681 72.7879
R6650 AVDD.n597 AVDD.n595 72.7879
R6651 AVDD.n602 AVDD.n600 72.7879
R6652 AVDD.n607 AVDD.n605 72.7879
R6653 AVDD.n613 AVDD.n610 72.7879
R6654 AVDD.n617 AVDD.n611 72.7879
R6655 AVDD.n622 AVDD.n620 72.7879
R6656 AVDD.n627 AVDD.n625 72.7879
R6657 AVDD.n632 AVDD.n630 72.7879
R6658 AVDD.n637 AVDD.n635 72.7879
R6659 AVDD.n642 AVDD.n640 72.7879
R6660 AVDD.n647 AVDD.n645 72.7879
R6661 AVDD.n652 AVDD.n650 72.7879
R6662 AVDD.n658 AVDD.n655 72.7879
R6663 AVDD.n662 AVDD.n656 72.7879
R6664 AVDD.n667 AVDD.n665 72.7879
R6665 AVDD.n672 AVDD.n670 72.7879
R6666 AVDD.n675 AVDD.n592 72.7879
R6667 AVDD.n3297 AVDD.n3296 56.1076
R6668 AVDD.n3297 AVDD.n14 56.1076
R6669 AVDD.n3297 AVDD.n15 56.1076
R6670 AVDD.n3297 AVDD.n16 56.1076
R6671 AVDD.n3297 AVDD.n17 56.1076
R6672 AVDD.n3297 AVDD.n18 56.1076
R6673 AVDD.n3297 AVDD.n19 56.1076
R6674 AVDD.n3297 AVDD.n20 56.1076
R6675 AVDD.n3297 AVDD.n21 56.1076
R6676 AVDD.n3297 AVDD.n22 56.1076
R6677 AVDD.n3297 AVDD.n23 56.1076
R6678 AVDD.n3297 AVDD.n24 56.1076
R6679 AVDD.n3297 AVDD.n25 56.1076
R6680 AVDD.n3297 AVDD.n26 56.1076
R6681 AVDD.n3297 AVDD.n27 56.1076
R6682 AVDD.n3297 AVDD.n28 56.1076
R6683 AVDD.n3297 AVDD.n29 56.1076
R6684 AVDD.n3297 AVDD.n30 56.1076
R6685 AVDD.n3297 AVDD.n31 56.1076
R6686 AVDD.n3297 AVDD.n32 56.1076
R6687 AVDD.n3297 AVDD.n33 56.1076
R6688 AVDD.n3297 AVDD.n34 56.1076
R6689 AVDD.n3297 AVDD.n35 56.1076
R6690 AVDD.n3297 AVDD.n36 56.1076
R6691 AVDD.n3297 AVDD.n37 56.1076
R6692 AVDD.n3297 AVDD.n38 56.1076
R6693 AVDD.n3297 AVDD.n39 56.1076
R6694 AVDD.n3297 AVDD.n40 56.1076
R6695 AVDD.n3297 AVDD.n41 56.1076
R6696 AVDD.n3297 AVDD.n43 56.1076
R6697 AVDD.n3297 AVDD.n44 56.1076
R6698 AVDD.n3297 AVDD.n45 56.1076
R6699 AVDD.n3297 AVDD.n46 56.1076
R6700 AVDD.n3297 AVDD.n47 56.1076
R6701 AVDD.n3297 AVDD.n48 56.1076
R6702 AVDD.n3297 AVDD.n49 56.1076
R6703 AVDD.n3297 AVDD.n50 56.1076
R6704 AVDD.n3297 AVDD.n51 56.1076
R6705 AVDD.n3297 AVDD.n52 56.1076
R6706 AVDD.n3297 AVDD.n53 56.1076
R6707 AVDD.n3297 AVDD.n54 56.1076
R6708 AVDD.n3297 AVDD.n55 56.1076
R6709 AVDD.n3297 AVDD.n56 56.1076
R6710 AVDD.n3297 AVDD.n57 56.1076
R6711 AVDD.n3297 AVDD.n58 56.1076
R6712 AVDD.n3297 AVDD.n59 56.1076
R6713 AVDD.n3297 AVDD.n60 56.1076
R6714 AVDD.n3297 AVDD.n61 56.1076
R6715 AVDD.n3297 AVDD.n63 56.1076
R6716 AVDD.n3297 AVDD.n64 56.1076
R6717 AVDD.n3297 AVDD.n65 56.1076
R6718 AVDD.n3297 AVDD.n66 56.1076
R6719 AVDD.n3297 AVDD.n67 56.1076
R6720 AVDD.n3297 AVDD.n68 56.1076
R6721 AVDD.n3297 AVDD.n69 56.1076
R6722 AVDD.n3297 AVDD.n70 56.1076
R6723 AVDD.n3297 AVDD.n71 56.1076
R6724 AVDD.n3297 AVDD.n72 56.1076
R6725 AVDD.n3297 AVDD.n73 56.1076
R6726 AVDD.n3297 AVDD.n74 56.1076
R6727 AVDD.n3297 AVDD.n75 56.1076
R6728 AVDD.n3297 AVDD.n76 56.1076
R6729 AVDD.n3297 AVDD.n77 56.1076
R6730 AVDD.n3297 AVDD.n78 56.1076
R6731 AVDD.n3298 AVDD.n3297 56.1076
R6732 AVDD.n3297 AVDD.n79 56.1076
R6733 AVDD.n3297 AVDD.n80 56.1076
R6734 AVDD.n3297 AVDD.n81 56.1076
R6735 AVDD.n3297 AVDD.n82 56.1076
R6736 AVDD.n3297 AVDD.n83 56.1076
R6737 AVDD.n3297 AVDD.n84 56.1076
R6738 AVDD.n3297 AVDD.n85 56.1076
R6739 AVDD.n3297 AVDD.n86 56.1076
R6740 AVDD.n3297 AVDD.n87 56.1076
R6741 AVDD.n3297 AVDD.n88 56.1076
R6742 AVDD.n3297 AVDD.n89 56.1076
R6743 AVDD.n3297 AVDD.n90 56.1076
R6744 AVDD.n3297 AVDD.n91 56.1076
R6745 AVDD.n491 AVDD.n200 56.1076
R6746 AVDD.n2843 AVDD.n200 56.1076
R6747 AVDD.n454 AVDD.n200 56.1076
R6748 AVDD.n2852 AVDD.n200 56.1076
R6749 AVDD.n445 AVDD.n200 56.1076
R6750 AVDD.n2862 AVDD.n200 56.1076
R6751 AVDD.n439 AVDD.n200 56.1076
R6752 AVDD.n2874 AVDD.n200 56.1076
R6753 AVDD.n424 AVDD.n200 56.1076
R6754 AVDD.n2884 AVDD.n200 56.1076
R6755 AVDD.n415 AVDD.n200 56.1076
R6756 AVDD.n2898 AVDD.n200 56.1076
R6757 AVDD.n407 AVDD.n200 56.1076
R6758 AVDD.n2908 AVDD.n200 56.1076
R6759 AVDD.n398 AVDD.n200 56.1076
R6760 AVDD.n2918 AVDD.n200 56.1076
R6761 AVDD.n376 AVDD.n200 56.1076
R6762 AVDD.n2928 AVDD.n200 56.1076
R6763 AVDD.n362 AVDD.n200 56.1076
R6764 AVDD.n2939 AVDD.n200 56.1076
R6765 AVDD.n356 AVDD.n200 56.1076
R6766 AVDD.n2948 AVDD.n200 56.1076
R6767 AVDD.n340 AVDD.n200 56.1076
R6768 AVDD.n2958 AVDD.n200 56.1076
R6769 AVDD.n332 AVDD.n200 56.1076
R6770 AVDD.n2968 AVDD.n200 56.1076
R6771 AVDD.n323 AVDD.n200 56.1076
R6772 AVDD.n2978 AVDD.n200 56.1076
R6773 AVDD.n317 AVDD.n200 56.1076
R6774 AVDD.n2990 AVDD.n200 56.1076
R6775 AVDD.n304 AVDD.n200 56.1076
R6776 AVDD.n3000 AVDD.n200 56.1076
R6777 AVDD.n292 AVDD.n200 56.1076
R6778 AVDD.n3014 AVDD.n200 56.1076
R6779 AVDD.n282 AVDD.n200 56.1076
R6780 AVDD.n3024 AVDD.n200 56.1076
R6781 AVDD.n275 AVDD.n200 56.1076
R6782 AVDD.n3036 AVDD.n200 56.1076
R6783 AVDD.n262 AVDD.n200 56.1076
R6784 AVDD.n3045 AVDD.n200 56.1076
R6785 AVDD.n252 AVDD.n200 56.1076
R6786 AVDD.n3059 AVDD.n200 56.1076
R6787 AVDD.n242 AVDD.n200 56.1076
R6788 AVDD.n3069 AVDD.n200 56.1076
R6789 AVDD.n235 AVDD.n200 56.1076
R6790 AVDD.n3081 AVDD.n200 56.1076
R6791 AVDD.n220 AVDD.n200 56.1076
R6792 AVDD.n3091 AVDD.n200 56.1076
R6793 AVDD.n213 AVDD.n200 56.1076
R6794 AVDD.n3101 AVDD.n200 56.1076
R6795 AVDD.n200 AVDD.n198 56.1076
R6796 AVDD.n1736 AVDD.n200 56.1076
R6797 AVDD.n1729 AVDD.n200 56.1076
R6798 AVDD.n1227 AVDD.n200 56.1076
R6799 AVDD.n1757 AVDD.n200 56.1076
R6800 AVDD.n1219 AVDD.n200 56.1076
R6801 AVDD.n1768 AVDD.n200 56.1076
R6802 AVDD.n1205 AVDD.n200 56.1076
R6803 AVDD.n1778 AVDD.n200 56.1076
R6804 AVDD.n1199 AVDD.n200 56.1076
R6805 AVDD.n1788 AVDD.n200 56.1076
R6806 AVDD.n1190 AVDD.n200 56.1076
R6807 AVDD.n1798 AVDD.n200 56.1076
R6808 AVDD.n1184 AVDD.n200 56.1076
R6809 AVDD.n1810 AVDD.n200 56.1076
R6810 AVDD.n1169 AVDD.n200 56.1076
R6811 AVDD.n1820 AVDD.n200 56.1076
R6812 AVDD.n1823 AVDD.n200 56.1076
R6813 AVDD.n1158 AVDD.n200 56.1076
R6814 AVDD.n1835 AVDD.n200 56.1076
R6815 AVDD.n1144 AVDD.n200 56.1076
R6816 AVDD.n1846 AVDD.n200 56.1076
R6817 AVDD.n549 AVDD.n200 56.1076
R6818 AVDD.n1856 AVDD.n200 56.1076
R6819 AVDD.n543 AVDD.n200 56.1076
R6820 AVDD.n1868 AVDD.n200 56.1076
R6821 AVDD.n530 AVDD.n200 56.1076
R6822 AVDD.n1877 AVDD.n200 56.1076
R6823 AVDD.n520 AVDD.n200 56.1076
R6824 AVDD.n1891 AVDD.n200 56.1076
R6825 AVDD.n845 AVDD.n776 56.1076
R6826 AVDD.n858 AVDD.n776 56.1076
R6827 AVDD.n839 AVDD.n776 56.1076
R6828 AVDD.n869 AVDD.n776 56.1076
R6829 AVDD.n832 AVDD.n776 56.1076
R6830 AVDD.n880 AVDD.n776 56.1076
R6831 AVDD.n889 AVDD.n776 56.1076
R6832 AVDD.n818 AVDD.n776 56.1076
R6833 AVDD.n898 AVDD.n776 56.1076
R6834 AVDD.n908 AVDD.n776 56.1076
R6835 AVDD.n805 AVDD.n776 56.1076
R6836 AVDD.n917 AVDD.n776 56.1076
R6837 AVDD.n928 AVDD.n776 56.1076
R6838 AVDD.n930 AVDD.n776 56.1076
R6839 AVDD.n939 AVDD.n776 56.1076
R6840 AVDD.n785 AVDD.n776 56.1076
R6841 AVDD.n964 AVDD.n776 56.1076
R6842 AVDD.n961 AVDD.n776 56.1076
R6843 AVDD.n951 AVDD.n776 56.1076
R6844 AVDD.n1137 AVDD.n1136 56.1076
R6845 AVDD.n1137 AVDD.n595 56.1076
R6846 AVDD.n1137 AVDD.n600 56.1076
R6847 AVDD.n1137 AVDD.n605 56.1076
R6848 AVDD.n1137 AVDD.n610 56.1076
R6849 AVDD.n1137 AVDD.n611 56.1076
R6850 AVDD.n1137 AVDD.n620 56.1076
R6851 AVDD.n1137 AVDD.n625 56.1076
R6852 AVDD.n1137 AVDD.n630 56.1076
R6853 AVDD.n1137 AVDD.n635 56.1076
R6854 AVDD.n1137 AVDD.n640 56.1076
R6855 AVDD.n1137 AVDD.n645 56.1076
R6856 AVDD.n1137 AVDD.n650 56.1076
R6857 AVDD.n1137 AVDD.n655 56.1076
R6858 AVDD.n1137 AVDD.n656 56.1076
R6859 AVDD.n1137 AVDD.n665 56.1076
R6860 AVDD.n1137 AVDD.n670 56.1076
R6861 AVDD.n1137 AVDD.n675 56.1076
R6862 AVDD.n1232 AVDD.n1230 56.0946
R6863 AVDD.n3124 AVDD.n185 56.0946
R6864 AVDD.n977 AVDD.n776 49.4282
R6865 AVDD.n1137 AVDD.n594 39.8722
R6866 AVDD.n1733 AVDD.n94 38.824
R6867 AVDD.n1734 AVDD.n1732 38.824
R6868 AVDD.n2362 AVDD.t110 28.5655
R6869 AVDD.n2362 AVDD.t53 28.5655
R6870 AVDD.n2604 AVDD.t288 28.5655
R6871 AVDD.n2604 AVDD.t389 28.5655
R6872 AVDD.n2603 AVDD.t196 28.5655
R6873 AVDD.t288 AVDD.n2603 28.5655
R6874 AVDD.n2579 AVDD.t254 28.5655
R6875 AVDD.n2579 AVDD.t196 28.5655
R6876 AVDD.n2538 AVDD.t208 28.5655
R6877 AVDD.n2538 AVDD.t189 28.5655
R6878 AVDD.n2537 AVDD.t397 28.5655
R6879 AVDD.t208 AVDD.n2537 28.5655
R6880 AVDD.n2476 AVDD.t406 28.5655
R6881 AVDD.n2476 AVDD.t397 28.5655
R6882 AVDD.n2475 AVDD.t299 28.5655
R6883 AVDD.t406 AVDD.n2475 28.5655
R6884 AVDD.n2474 AVDD.t217 28.5655
R6885 AVDD.t299 AVDD.n2474 28.5655
R6886 AVDD.n2427 AVDD.t212 28.5655
R6887 AVDD.n2427 AVDD.t294 28.5655
R6888 AVDD.n2426 AVDD.t222 28.5655
R6889 AVDD.t212 AVDD.n2426 28.5655
R6890 AVDD.t411 AVDD.n2386 28.5655
R6891 AVDD.n2386 AVDD.t222 28.5655
R6892 AVDD.t335 AVDD.n1883 28.5655
R6893 AVDD.n1883 AVDD.t324 28.5655
R6894 AVDD.t200 AVDD.n537 28.5655
R6895 AVDD.n537 AVDD.t186 28.5655
R6896 AVDD.t379 AVDD.n1152 28.5655
R6897 AVDD.n1152 AVDD.t361 28.5655
R6898 AVDD.t147 AVDD.n1178 28.5655
R6899 AVDD.n1178 AVDD.t135 28.5655
R6900 AVDD.t310 AVDD.n1212 28.5655
R6901 AVDD.n1212 AVDD.t307 28.5655
R6902 AVDD.t165 AVDD.n1235 28.5655
R6903 AVDD.n1235 AVDD.t156 28.5655
R6904 AVDD.t181 AVDD.n206 28.5655
R6905 AVDD.n206 AVDD.t175 28.5655
R6906 AVDD.t343 AVDD.n229 28.5655
R6907 AVDD.n229 AVDD.t337 28.5655
R6908 AVDD.t169 AVDD.n3051 28.5655
R6909 AVDD.n3051 AVDD.t159 28.5655
R6910 AVDD.t330 AVDD.n269 28.5655
R6911 AVDD.n269 AVDD.t321 28.5655
R6912 AVDD.t284 AVDD.n3006 28.5655
R6913 AVDD.n3006 AVDD.t214 28.5655
R6914 AVDD.t418 AVDD.n311 28.5655
R6915 AVDD.n311 AVDD.t332 28.5655
R6916 AVDD.t171 AVDD.n347 28.5655
R6917 AVDD.n347 AVDD.t162 28.5655
R6918 AVDD.t232 AVDD.n369 28.5655
R6919 AVDD.n369 AVDD.t315 28.5655
R6920 AVDD.t142 AVDD.n2890 28.5655
R6921 AVDD.n2890 AVDD.t244 28.5655
R6922 AVDD.t282 AVDD.n433 28.5655
R6923 AVDD.n433 AVDD.t367 28.5655
R6924 AVDD.t269 AVDD.n460 28.5655
R6925 AVDD.n460 AVDD.t353 28.5655
R6926 AVDD.n1069 AVDD.t264 28.5655
R6927 AVDD.n1069 AVDD.t327 28.5655
R6928 AVDD.n1068 AVDD.t273 28.5655
R6929 AVDD.t264 AVDD.n1068 28.5655
R6930 AVDD.t167 AVDD.n1009 28.5655
R6931 AVDD.n1009 AVDD.t258 28.5655
R6932 AVDD.n1010 AVDD.t173 28.5655
R6933 AVDD.n1010 AVDD.t167 28.5655
R6934 AVDD.t236 AVDD.n103 28.5655
R6935 AVDD.n103 AVDD.t227 28.5655
R6936 AVDD.t416 AVDD.n116 28.5655
R6937 AVDD.n116 AVDD.t408 28.5655
R6938 AVDD.t277 AVDD.n133 28.5655
R6939 AVDD.n133 AVDD.t266 28.5655
R6940 AVDD.t345 AVDD.n151 28.5655
R6941 AVDD.n151 AVDD.t340 28.5655
R6942 AVDD.t210 AVDD.n3153 28.5655
R6943 AVDD.n3153 AVDD.t205 28.5655
R6944 AVDD.t381 AVDD.n182 28.5655
R6945 AVDD.n182 AVDD.t364 28.5655
R6946 AVDD.t404 AVDD.n1339 28.5655
R6947 AVDD.n1339 AVDD.t399 28.5655
R6948 AVDD.t252 AVDD.n1324 28.5655
R6949 AVDD.n1324 AVDD.t241 28.5655
R6950 AVDD.t387 AVDD.n1683 28.5655
R6951 AVDD.n1683 AVDD.t373 28.5655
R6952 AVDD.t230 AVDD.n1405 28.5655
R6953 AVDD.n1405 AVDD.t219 28.5655
R6954 AVDD.t271 AVDD.n1628 28.5655
R6955 AVDD.n1628 AVDD.t193 28.5655
R6956 AVDD.t402 AVDD.n1456 28.5655
R6957 AVDD.n1456 AVDD.t312 28.5655
R6958 AVDD.t392 AVDD.n1561 28.5655
R6959 AVDD.n1561 AVDD.t376 28.5655
R6960 AVDD.t234 AVDD.n1510 28.5655
R6961 AVDD.n1510 AVDD.t318 28.5655
R6962 AVDD.t145 AVDD.n2248 28.5655
R6963 AVDD.n2248 AVDD.t247 28.5655
R6964 AVDD.t286 AVDD.n2282 28.5655
R6965 AVDD.n2282 AVDD.t370 28.5655
R6966 AVDD.t275 AVDD.n2216 28.5655
R6967 AVDD.n2216 AVDD.t356 28.5655
R6968 AVDD.n2140 AVDD.t250 28.5655
R6969 AVDD.n2140 AVDD.t238 28.5655
R6970 AVDD.n2139 AVDD.t256 28.5655
R6971 AVDD.t250 AVDD.n2139 28.5655
R6972 AVDD.n2138 AVDD.t383 28.5655
R6973 AVDD.t256 AVDD.n2138 28.5655
R6974 AVDD.n2071 AVDD.t385 28.5655
R6975 AVDD.n2071 AVDD.t138 28.5655
R6976 AVDD.n2070 AVDD.t359 28.5655
R6977 AVDD.t385 AVDD.n2070 28.5655
R6978 AVDD.n2069 AVDD.t290 28.5655
R6979 AVDD.t359 AVDD.n2069 28.5655
R6980 AVDD.n2068 AVDD.t292 28.5655
R6981 AVDD.t290 AVDD.n2068 28.5655
R6982 AVDD.n2065 AVDD.t297 28.5655
R6983 AVDD.t292 AVDD.n2065 28.5655
R6984 AVDD.n1974 AVDD.t198 28.5655
R6985 AVDD.n1974 AVDD.t178 28.5655
R6986 AVDD.n1973 AVDD.t128 28.5655
R6987 AVDD.t198 AVDD.n1973 28.5655
R6988 AVDD.n1970 AVDD.t420 28.5655
R6989 AVDD.t128 AVDD.n1970 28.5655
R6990 AVDD.n1261 AVDD.t113 28.5655
R6991 AVDD.n1261 AVDD.t123 28.5655
R6992 AVDD.n1260 AVDD.t54 28.5655
R6993 AVDD.n1260 AVDD.t64 28.5655
R6994 AVDD.n1286 AVDD.t86 28.5655
R6995 AVDD.n1286 AVDD.t94 28.5655
R6996 AVDD.n1285 AVDD.t34 28.5655
R6997 AVDD.n1285 AVDD.t45 28.5655
R6998 AVDD.n1245 AVDD.t48 28.5655
R6999 AVDD.n1245 AVDD.t56 28.5655
R7000 AVDD.n1244 AVDD.t80 28.5655
R7001 AVDD.n1244 AVDD.t85 28.5655
R7002 AVDD.n1312 AVDD.t111 28.5655
R7003 AVDD.n1312 AVDD.t120 28.5655
R7004 AVDD.n1311 AVDD.t33 28.5655
R7005 AVDD.n1311 AVDD.t42 28.5655
R7006 AVDD.n1423 AVDD.t101 28.5655
R7007 AVDD.n1423 AVDD.t63 28.5655
R7008 AVDD.n1422 AVDD.t97 28.5655
R7009 AVDD.n1422 AVDD.t105 28.5655
R7010 AVDD.n1477 AVDD.t49 28.5655
R7011 AVDD.n1477 AVDD.t58 28.5655
R7012 AVDD.n1476 AVDD.t115 28.5655
R7013 AVDD.n1476 AVDD.t74 28.5655
R7014 AVDD.n387 AVDD.t71 28.5655
R7015 AVDD.n387 AVDD.t114 28.5655
R7016 AVDD.n386 AVDD.t91 28.5655
R7017 AVDD.n386 AVDD.t36 28.5655
R7018 AVDD.n1746 AVDD.n200 28.0408
R7019 AVDD.n1106 AVDD.n684 27.3755
R7020 AVDD.n3089 AVDD.n214 25.6005
R7021 AVDD.n260 AVDD.n256 25.6005
R7022 AVDD.n2988 AVDD.n305 25.6005
R7023 AVDD.n354 AVDD.n344 25.6005
R7024 AVDD.n2896 AVDD.n408 25.6005
R7025 AVDD.n452 AVDD.n449 25.6005
R7026 AVDD.n1362 AVDD.n1359 25.6005
R7027 AVDD.n1669 AVDD.n1666 25.6005
R7028 AVDD.n1451 AVDD.n1447 25.6005
R7029 AVDD.n1502 AVDD.n1498 25.6005
R7030 AVDD.n2244 AVDD.n2232 25.6005
R7031 AVDD.n2317 AVDD.n2314 25.6005
R7032 AVDD.n2409 AVDD.n2401 25.6005
R7033 AVDD.n2463 AVDD.n2458 25.6005
R7034 AVDD.n2558 AVDD.n2555 25.6005
R7035 AVDD.n2624 AVDD.n2621 25.6005
R7036 AVDD.n528 AVDD.n524 25.6005
R7037 AVDD.n1825 AVDD.n1157 25.6005
R7038 AVDD.n1776 AVDD.n1200 25.6005
R7039 AVDD.n2404 AVDD.n1949 25.6005
R7040 AVDD.n2465 AVDD.n2013 25.6005
R7041 AVDD.n2088 AVDD.n2082 25.6005
R7042 AVDD.n2157 AVDD.n2151 25.6005
R7043 AVDD.n3276 AVDD.n3273 25.6005
R7044 AVDD.n3221 AVDD.n3218 25.6005
R7045 AVDD.n3169 AVDD.n3166 25.6005
R7046 AVDD.n932 AVDD.n796 25.6005
R7047 AVDD.n837 AVDD.n833 25.6005
R7048 AVDD.n1058 AVDD.n1057 25.6005
R7049 AVDD.n616 AVDD.n615 25.6005
R7050 AVDD.n661 AVDD.n660 25.6005
R7051 AVDD.n1049 AVDD.n1048 25.6005
R7052 AVDD.n1056 AVDD.n1051 25.224
R7053 AVDD.n1040 AVDD.n745 25.224
R7054 AVDD.n3094 AVDD.n212 24.8476
R7055 AVDD.n3088 AVDD.n216 24.8476
R7056 AVDD.n3043 AVDD.n3042 24.8476
R7057 AVDD.n3039 AVDD.n3038 24.8476
R7058 AVDD.n2993 AVDD.n302 24.8476
R7059 AVDD.n2987 AVDD.n307 24.8476
R7060 AVDD.n2946 AVDD.n2945 24.8476
R7061 AVDD.n2942 AVDD.n2941 24.8476
R7062 AVDD.n2901 AVDD.n406 24.8476
R7063 AVDD.n2895 AVDD.n410 24.8476
R7064 AVDD.n2850 AVDD.n2849 24.8476
R7065 AVDD.n2846 AVDD.n2845 24.8476
R7066 AVDD.n1358 AVDD.n1330 24.8476
R7067 AVDD.n1366 AVDD.n1363 24.8476
R7068 AVDD.n1673 AVDD.n1670 24.8476
R7069 AVDD.n1665 AVDD.n1399 24.8476
R7070 AVDD.n1614 AVDD.n1612 24.8476
R7071 AVDD.n1609 AVDD.n1608 24.8476
R7072 AVDD.n1558 AVDD.n1555 24.8476
R7073 AVDD.n1552 AVDD.n1551 24.8476
R7074 AVDD.n2245 AVDD.n2241 24.8476
R7075 AVDD.n2256 AVDD.n2253 24.8476
R7076 AVDD.n2313 AVDD.n2219 24.8476
R7077 AVDD.n2319 AVDD.n2318 24.8476
R7078 AVDD.n2410 AVDD.n2399 24.8476
R7079 AVDD.n2400 AVDD.n2381 24.8476
R7080 AVDD.n2509 AVDD.n2508 24.8476
R7081 AVDD.n2470 AVDD.n2461 24.8476
R7082 AVDD.n2554 AVDD.n2357 24.8476
R7083 AVDD.n2559 AVDD.n2355 24.8476
R7084 AVDD.n2620 AVDD.n2338 24.8476
R7085 AVDD.n2625 AVDD.n2211 24.8476
R7086 AVDD.n1875 AVDD.n1874 24.8476
R7087 AVDD.n1871 AVDD.n1870 24.8476
R7088 AVDD.n1826 AVDD.n1156 24.8476
R7089 AVDD.n1161 AVDD.n1160 24.8476
R7090 AVDD.n1781 AVDD.n1198 24.8476
R7091 AVDD.n1775 AVDD.n1202 24.8476
R7092 AVDD.n2817 AVDD.n2816 24.8476
R7093 AVDD.n2403 AVDD.n1957 24.8476
R7094 AVDD.n2766 AVDD.n2765 24.8476
R7095 AVDD.n2464 AVDD.n2021 24.8476
R7096 AVDD.n2714 AVDD.n2713 24.8476
R7097 AVDD.n2709 AVDD.n2708 24.8476
R7098 AVDD.n2663 AVDD.n2662 24.8476
R7099 AVDD.n2658 AVDD.n2657 24.8476
R7100 AVDD.n3280 AVDD.n3277 24.8476
R7101 AVDD.n3272 AVDD.n110 24.8476
R7102 AVDD.n3222 AVDD.n139 24.8476
R7103 AVDD.n3217 AVDD.n3216 24.8476
R7104 AVDD.n3173 AVDD.n3170 24.8476
R7105 AVDD.n3165 AVDD.n166 24.8476
R7106 AVDD.n933 AVDD.n793 24.8476
R7107 AVDD.n926 AVDD.n798 24.8476
R7108 AVDD.n878 AVDD.n877 24.8476
R7109 AVDD.n872 AVDD.n871 24.8476
R7110 AVDD.n612 AVDD.n568 24.8476
R7111 AVDD.n618 AVDD.n583 24.8476
R7112 AVDD.n657 AVDD.n573 24.8476
R7113 AVDD.n663 AVDD.n587 24.8476
R7114 AVDD.n303 AVDD.n295 24.7064
R7115 AVDD.n294 AVDD.n93 24.7064
R7116 AVDD.n1076 AVDD.n732 24.4711
R7117 AVDD.n1047 AVDD.n726 24.4711
R7118 AVDD.n1064 AVDD.n738 23.7181
R7119 AVDD.n1041 AVDD.n1039 23.7181
R7120 AVDD.n3095 AVDD.n203 23.3417
R7121 AVDD.n3085 AVDD.n3084 23.3417
R7122 AVDD.n255 AVDD.n253 23.3417
R7123 AVDD.n3034 AVDD.n261 23.3417
R7124 AVDD.n2994 AVDD.n297 23.3417
R7125 AVDD.n315 AVDD.n314 23.3417
R7126 AVDD.n343 AVDD.n341 23.3417
R7127 AVDD.n2937 AVDD.n355 23.3417
R7128 AVDD.n2902 AVDD.n402 23.3417
R7129 AVDD.n2888 AVDD.n2887 23.3417
R7130 AVDD.n448 AVDD.n446 23.3417
R7131 AVDD.n2841 AVDD.n453 23.3417
R7132 AVDD.n1354 AVDD.n1353 23.3417
R7133 AVDD.n1367 AVDD.n1328 23.3417
R7134 AVDD.n1674 AVDD.n1397 23.3417
R7135 AVDD.n1661 AVDD.n1660 23.3417
R7136 AVDD.n1615 AVDD.n1446 23.3417
R7137 AVDD.n1605 AVDD.n1452 23.3417
R7138 AVDD.n1559 AVDD.n1495 23.3417
R7139 AVDD.n1548 AVDD.n1503 23.3417
R7140 AVDD.n2238 AVDD.n2234 23.3417
R7141 AVDD.n2257 AVDD.n2230 23.3417
R7142 AVDD.n2310 AVDD.n2309 23.3417
R7143 AVDD.n2330 AVDD.n2329 23.3417
R7144 AVDD.n2398 AVDD.n2384 23.3417
R7145 AVDD.n2417 AVDD.n2416 23.3417
R7146 AVDD.n2510 AVDD.n2457 23.3417
R7147 AVDD.n2502 AVDD.n2501 23.3417
R7148 AVDD.n2547 AVDD.n2546 23.3417
R7149 AVDD.n2563 AVDD.n2562 23.3417
R7150 AVDD.n2613 AVDD.n2612 23.3417
R7151 AVDD.n2634 AVDD.n2633 23.3417
R7152 AVDD.n523 AVDD.n521 23.3417
R7153 AVDD.n1866 AVDD.n529 23.3417
R7154 AVDD.n1155 AVDD.n1148 23.3417
R7155 AVDD.n1818 AVDD.n1163 23.3417
R7156 AVDD.n1782 AVDD.n1194 23.3417
R7157 AVDD.n1772 AVDD.n1771 23.3417
R7158 AVDD.n1948 AVDD.n1947 23.3417
R7159 AVDD.n2810 AVDD.n2809 23.3417
R7160 AVDD.n2012 AVDD.n2011 23.3417
R7161 AVDD.n2759 AVDD.n2758 23.3417
R7162 AVDD.n2081 AVDD.n2080 23.3417
R7163 AVDD.n2098 AVDD.n2089 23.3417
R7164 AVDD.n2150 AVDD.n2149 23.3417
R7165 AVDD.n2167 AVDD.n2158 23.3417
R7166 AVDD.n3281 AVDD.n108 23.3417
R7167 AVDD.n3268 AVDD.n3267 23.3417
R7168 AVDD.n136 AVDD.n129 23.3417
R7169 AVDD.n3213 AVDD.n140 23.3417
R7170 AVDD.n3174 AVDD.n162 23.3417
R7171 AVDD.n3162 AVDD.n3161 23.3417
R7172 AVDD.n937 AVDD.n936 23.3417
R7173 AVDD.n925 AVDD.n799 23.3417
R7174 AVDD.n882 AVDD.n831 23.3417
R7175 AVDD.n865 AVDD.n838 23.3417
R7176 AVDD.n608 AVDD.n578 23.3417
R7177 AVDD.n621 AVDD.n562 23.3417
R7178 AVDD.n653 AVDD.n572 23.3417
R7179 AVDD.n666 AVDD.n558 23.3417
R7180 AVDD.n1075 AVDD.n733 22.9652
R7181 AVDD.n1082 AVDD.n1081 22.9652
R7182 AVDD.n1885 AVDD.n516 22.5538
R7183 AVDD.n517 AVDD.n516 22.5538
R7184 AVDD.n1884 AVDD.n516 22.5538
R7185 AVDD.n1863 AVDD.n1862 22.5538
R7186 AVDD.n1863 AVDD.n535 22.5538
R7187 AVDD.n1863 AVDD.n538 22.5538
R7188 AVDD.n1830 AVDD.n1829 22.5538
R7189 AVDD.n1830 AVDD.n1150 22.5538
R7190 AVDD.n1830 AVDD.n1153 22.5538
R7191 AVDD.n1805 AVDD.n1804 22.5538
R7192 AVDD.n1805 AVDD.n1176 22.5538
R7193 AVDD.n1805 AVDD.n1179 22.5538
R7194 AVDD.n1214 AVDD.n1203 22.5538
R7195 AVDD.n1211 AVDD.n1203 22.5538
R7196 AVDD.n1213 AVDD.n1203 22.5538
R7197 AVDD.n1238 AVDD.n1237 22.5538
R7198 AVDD.n1237 AVDD.n1234 22.5538
R7199 AVDD.n1237 AVDD.n1236 22.5538
R7200 AVDD.n209 AVDD.n208 22.5538
R7201 AVDD.n208 AVDD.n205 22.5538
R7202 AVDD.n208 AVDD.n207 22.5538
R7203 AVDD.n3076 AVDD.n3075 22.5538
R7204 AVDD.n3076 AVDD.n227 22.5538
R7205 AVDD.n3076 AVDD.n230 22.5538
R7206 AVDD.n3053 AVDD.n248 22.5538
R7207 AVDD.n249 AVDD.n248 22.5538
R7208 AVDD.n3052 AVDD.n248 22.5538
R7209 AVDD.n3031 AVDD.n3030 22.5538
R7210 AVDD.n3031 AVDD.n267 22.5538
R7211 AVDD.n3031 AVDD.n270 22.5538
R7212 AVDD.n3008 AVDD.n288 22.5538
R7213 AVDD.n289 AVDD.n288 22.5538
R7214 AVDD.n3007 AVDD.n288 22.5538
R7215 AVDD.n2985 AVDD.n2984 22.5538
R7216 AVDD.n2985 AVDD.n309 22.5538
R7217 AVDD.n2985 AVDD.n312 22.5538
R7218 AVDD.n349 AVDD.n338 22.5538
R7219 AVDD.n346 AVDD.n338 22.5538
R7220 AVDD.n348 AVDD.n338 22.5538
R7221 AVDD.n372 AVDD.n371 22.5538
R7222 AVDD.n371 AVDD.n368 22.5538
R7223 AVDD.n371 AVDD.n370 22.5538
R7224 AVDD.n2892 AVDD.n411 22.5538
R7225 AVDD.n412 AVDD.n411 22.5538
R7226 AVDD.n2891 AVDD.n411 22.5538
R7227 AVDD.n2869 AVDD.n2868 22.5538
R7228 AVDD.n2869 AVDD.n431 22.5538
R7229 AVDD.n2869 AVDD.n434 22.5538
R7230 AVDD.n462 AVDD.n458 22.5538
R7231 AVDD.n459 AVDD.n458 22.5538
R7232 AVDD.n461 AVDD.n458 22.5538
R7233 AVDD.n944 AVDD.n787 22.5538
R7234 AVDD.n788 AVDD.n787 22.5538
R7235 AVDD.n922 AVDD.n801 22.5538
R7236 AVDD.n802 AVDD.n801 22.5538
R7237 AVDD.n814 AVDD.n807 22.5538
R7238 AVDD.n813 AVDD.n807 22.5538
R7239 AVDD.n828 AVDD.n821 22.5538
R7240 AVDD.n827 AVDD.n821 22.5538
R7241 AVDD.n874 AVDD.n834 22.5538
R7242 AVDD.n835 AVDD.n834 22.5538
R7243 AVDD.n853 AVDD.n852 22.5538
R7244 AVDD.n853 AVDD.n849 22.5538
R7245 AVDD.n3291 AVDD.n3290 22.5538
R7246 AVDD.n3291 AVDD.n101 22.5538
R7247 AVDD.n3291 AVDD.n104 22.5538
R7248 AVDD.n119 AVDD.n118 22.5538
R7249 AVDD.n118 AVDD.n115 22.5538
R7250 AVDD.n118 AVDD.n117 22.5538
R7251 AVDD.n3226 AVDD.n3225 22.5538
R7252 AVDD.n3226 AVDD.n131 22.5538
R7253 AVDD.n3226 AVDD.n134 22.5538
R7254 AVDD.n3198 AVDD.n3197 22.5538
R7255 AVDD.n3198 AVDD.n149 22.5538
R7256 AVDD.n3198 AVDD.n152 22.5538
R7257 AVDD.n3155 AVDD.n167 22.5538
R7258 AVDD.n169 AVDD.n167 22.5538
R7259 AVDD.n3154 AVDD.n167 22.5538
R7260 AVDD.n3128 AVDD.n3127 22.5538
R7261 AVDD.n3128 AVDD.n180 22.5538
R7262 AVDD.n3128 AVDD.n183 22.5538
R7263 AVDD.n1343 AVDD.n1342 22.5538
R7264 AVDD.n1343 AVDD.n1337 22.5538
R7265 AVDD.n1343 AVDD.n1340 22.5538
R7266 AVDD.n1383 AVDD.n1382 22.5538
R7267 AVDD.n1382 AVDD.n1323 22.5538
R7268 AVDD.n1382 AVDD.n1325 22.5538
R7269 AVDD.n1685 AVDD.n1393 22.5538
R7270 AVDD.n1395 AVDD.n1393 22.5538
R7271 AVDD.n1684 AVDD.n1393 22.5538
R7272 AVDD.n1408 AVDD.n1407 22.5538
R7273 AVDD.n1407 AVDD.n1404 22.5538
R7274 AVDD.n1407 AVDD.n1406 22.5538
R7275 AVDD.n1630 AVDD.n1440 22.5538
R7276 AVDD.n1441 AVDD.n1440 22.5538
R7277 AVDD.n1629 AVDD.n1440 22.5538
R7278 AVDD.n1458 AVDD.n1448 22.5538
R7279 AVDD.n1455 AVDD.n1448 22.5538
R7280 AVDD.n1457 AVDD.n1448 22.5538
R7281 AVDD.n1563 AVDD.n1494 22.5538
R7282 AVDD.n1496 AVDD.n1494 22.5538
R7283 AVDD.n1562 AVDD.n1494 22.5538
R7284 AVDD.n1513 AVDD.n1512 22.5538
R7285 AVDD.n1512 AVDD.n1509 22.5538
R7286 AVDD.n1512 AVDD.n1511 22.5538
R7287 AVDD.n2251 AVDD.n2250 22.5538
R7288 AVDD.n2251 AVDD.n2247 22.5538
R7289 AVDD.n2251 AVDD.n2249 22.5538
R7290 AVDD.n2286 AVDD.n2285 22.5538
R7291 AVDD.n2286 AVDD.n2280 22.5538
R7292 AVDD.n2286 AVDD.n2283 22.5538
R7293 AVDD.n2333 AVDD.n2332 22.5538
R7294 AVDD.n2332 AVDD.n2214 22.5538
R7295 AVDD.n2332 AVDD.n2217 22.5538
R7296 AVDD.n1886 AVDD.n1885 22.5534
R7297 AVDD.n1886 AVDD.n517 22.5534
R7298 AVDD.n1886 AVDD.n1884 22.5534
R7299 AVDD.n1862 AVDD.n1861 22.5534
R7300 AVDD.n1861 AVDD.n535 22.5534
R7301 AVDD.n1861 AVDD.n538 22.5534
R7302 AVDD.n1829 AVDD.n1828 22.5534
R7303 AVDD.n1828 AVDD.n1150 22.5534
R7304 AVDD.n1828 AVDD.n1153 22.5534
R7305 AVDD.n1804 AVDD.n1803 22.5534
R7306 AVDD.n1803 AVDD.n1176 22.5534
R7307 AVDD.n1803 AVDD.n1179 22.5534
R7308 AVDD.n1215 AVDD.n1214 22.5534
R7309 AVDD.n1215 AVDD.n1211 22.5534
R7310 AVDD.n1215 AVDD.n1213 22.5534
R7311 AVDD.n1239 AVDD.n1238 22.5534
R7312 AVDD.n1239 AVDD.n1234 22.5534
R7313 AVDD.n1239 AVDD.n1236 22.5534
R7314 AVDD.n210 AVDD.n209 22.5534
R7315 AVDD.n210 AVDD.n205 22.5534
R7316 AVDD.n210 AVDD.n207 22.5534
R7317 AVDD.n3075 AVDD.n3074 22.5534
R7318 AVDD.n3074 AVDD.n227 22.5534
R7319 AVDD.n3074 AVDD.n230 22.5534
R7320 AVDD.n3054 AVDD.n3053 22.5534
R7321 AVDD.n3054 AVDD.n249 22.5534
R7322 AVDD.n3054 AVDD.n3052 22.5534
R7323 AVDD.n3030 AVDD.n3029 22.5534
R7324 AVDD.n3029 AVDD.n267 22.5534
R7325 AVDD.n3029 AVDD.n270 22.5534
R7326 AVDD.n3009 AVDD.n3008 22.5534
R7327 AVDD.n3009 AVDD.n289 22.5534
R7328 AVDD.n3009 AVDD.n3007 22.5534
R7329 AVDD.n2984 AVDD.n2983 22.5534
R7330 AVDD.n2983 AVDD.n309 22.5534
R7331 AVDD.n2983 AVDD.n312 22.5534
R7332 AVDD.n350 AVDD.n349 22.5534
R7333 AVDD.n350 AVDD.n346 22.5534
R7334 AVDD.n350 AVDD.n348 22.5534
R7335 AVDD.n373 AVDD.n372 22.5534
R7336 AVDD.n373 AVDD.n368 22.5534
R7337 AVDD.n373 AVDD.n370 22.5534
R7338 AVDD.n2893 AVDD.n2892 22.5534
R7339 AVDD.n2893 AVDD.n412 22.5534
R7340 AVDD.n2893 AVDD.n2891 22.5534
R7341 AVDD.n2868 AVDD.n2867 22.5534
R7342 AVDD.n2867 AVDD.n431 22.5534
R7343 AVDD.n2867 AVDD.n434 22.5534
R7344 AVDD.n463 AVDD.n462 22.5534
R7345 AVDD.n463 AVDD.n459 22.5534
R7346 AVDD.n463 AVDD.n461 22.5534
R7347 AVDD.n945 AVDD.n944 22.5534
R7348 AVDD.n945 AVDD.n788 22.5534
R7349 AVDD.n923 AVDD.n922 22.5534
R7350 AVDD.n923 AVDD.n802 22.5534
R7351 AVDD.n815 AVDD.n814 22.5534
R7352 AVDD.n815 AVDD.n813 22.5534
R7353 AVDD.n829 AVDD.n828 22.5534
R7354 AVDD.n829 AVDD.n827 22.5534
R7355 AVDD.n875 AVDD.n874 22.5534
R7356 AVDD.n875 AVDD.n835 22.5534
R7357 AVDD.n852 AVDD.n773 22.5534
R7358 AVDD.n849 AVDD.n773 22.5534
R7359 AVDD.n3290 AVDD.n3289 22.5534
R7360 AVDD.n3289 AVDD.n101 22.5534
R7361 AVDD.n3289 AVDD.n104 22.5534
R7362 AVDD.n120 AVDD.n119 22.5534
R7363 AVDD.n120 AVDD.n115 22.5534
R7364 AVDD.n120 AVDD.n117 22.5534
R7365 AVDD.n3225 AVDD.n3224 22.5534
R7366 AVDD.n3224 AVDD.n131 22.5534
R7367 AVDD.n3224 AVDD.n134 22.5534
R7368 AVDD.n3197 AVDD.n3196 22.5534
R7369 AVDD.n3196 AVDD.n149 22.5534
R7370 AVDD.n3196 AVDD.n152 22.5534
R7371 AVDD.n3156 AVDD.n3155 22.5534
R7372 AVDD.n3156 AVDD.n169 22.5534
R7373 AVDD.n3156 AVDD.n3154 22.5534
R7374 AVDD.n3127 AVDD.n3126 22.5534
R7375 AVDD.n3126 AVDD.n180 22.5534
R7376 AVDD.n3126 AVDD.n183 22.5534
R7377 AVDD.n1342 AVDD.n1341 22.5534
R7378 AVDD.n1341 AVDD.n1337 22.5534
R7379 AVDD.n1341 AVDD.n1340 22.5534
R7380 AVDD.n1384 AVDD.n1383 22.5534
R7381 AVDD.n1384 AVDD.n1323 22.5534
R7382 AVDD.n1384 AVDD.n1325 22.5534
R7383 AVDD.n1686 AVDD.n1685 22.5534
R7384 AVDD.n1686 AVDD.n1395 22.5534
R7385 AVDD.n1686 AVDD.n1684 22.5534
R7386 AVDD.n1409 AVDD.n1408 22.5534
R7387 AVDD.n1409 AVDD.n1404 22.5534
R7388 AVDD.n1409 AVDD.n1406 22.5534
R7389 AVDD.n1631 AVDD.n1630 22.5534
R7390 AVDD.n1631 AVDD.n1441 22.5534
R7391 AVDD.n1631 AVDD.n1629 22.5534
R7392 AVDD.n1459 AVDD.n1458 22.5534
R7393 AVDD.n1459 AVDD.n1455 22.5534
R7394 AVDD.n1459 AVDD.n1457 22.5534
R7395 AVDD.n1564 AVDD.n1563 22.5534
R7396 AVDD.n1564 AVDD.n1496 22.5534
R7397 AVDD.n1564 AVDD.n1562 22.5534
R7398 AVDD.n1514 AVDD.n1513 22.5534
R7399 AVDD.n1514 AVDD.n1509 22.5534
R7400 AVDD.n1514 AVDD.n1511 22.5534
R7401 AVDD.n2250 AVDD.n2231 22.5534
R7402 AVDD.n2247 AVDD.n2231 22.5534
R7403 AVDD.n2249 AVDD.n2231 22.5534
R7404 AVDD.n2285 AVDD.n2284 22.5534
R7405 AVDD.n2284 AVDD.n2280 22.5534
R7406 AVDD.n2284 AVDD.n2283 22.5534
R7407 AVDD.n2334 AVDD.n2333 22.5534
R7408 AVDD.n2334 AVDD.n2214 22.5534
R7409 AVDD.n2334 AVDD.n2217 22.5534
R7410 AVDD.n977 AVDD.n777 22.4077
R7411 AVDD.n986 AVDD.n763 22.4077
R7412 AVDD.n999 AVDD.n763 22.4077
R7413 AVDD.n999 AVDD.n756 22.4077
R7414 AVDD.n1021 AVDD.n756 22.4077
R7415 AVDD.n1021 AVDD.n1020 22.4077
R7416 AVDD.n1034 AVDD.n741 22.4077
R7417 AVDD.n1062 AVDD.n741 22.4077
R7418 AVDD.n1062 AVDD.n1061 22.4077
R7419 AVDD.n1060 AVDD.n730 22.4077
R7420 AVDD.n1078 AVDD.n730 22.4077
R7421 AVDD.n1079 AVDD.n1078 22.4077
R7422 AVDD.n1094 AVDD.n1093 22.4077
R7423 AVDD.n1093 AVDD.n708 22.4077
R7424 AVDD.n1111 AVDD.n708 22.4077
R7425 AVDD.n1111 AVDD.n689 22.4077
R7426 AVDD.n1122 AVDD.n689 22.4077
R7427 AVDD.n1123 AVDD.n1122 22.4077
R7428 AVDD.n1126 AVDD.n594 22.4077
R7429 AVDD.n1065 AVDD.n737 22.2123
R7430 AVDD.n1038 AVDD.n1037 22.2123
R7431 AVDD.n2617 AVDD.n2616 21.9522
R7432 AVDD.n2618 AVDD.n2617 21.9522
R7433 AVDD.n2345 AVDD.n2344 21.9522
R7434 AVDD.n2344 AVDD.n2342 21.9522
R7435 AVDD.n2589 AVDD.n2588 21.9522
R7436 AVDD.n2590 AVDD.n2589 21.9522
R7437 AVDD.n2573 AVDD.n2572 21.9522
R7438 AVDD.n2572 AVDD.n2349 21.9522
R7439 AVDD.n2551 AVDD.n2550 21.9522
R7440 AVDD.n2552 AVDD.n2551 21.9522
R7441 AVDD.n2530 AVDD.n2529 21.9522
R7442 AVDD.n2529 AVDD.n2361 21.9522
R7443 AVDD.n2483 AVDD.n2482 21.9522
R7444 AVDD.n2482 AVDD.n2367 21.9522
R7445 AVDD.n2496 AVDD.n2495 21.9522
R7446 AVDD.n2495 AVDD.n2494 21.9522
R7447 AVDD.n2506 AVDD.n2505 21.9522
R7448 AVDD.n2505 AVDD.n2504 21.9522
R7449 AVDD.n2514 AVDD.n2513 21.9522
R7450 AVDD.n2513 AVDD.n2512 21.9522
R7451 AVDD.n2437 AVDD.n2436 21.9522
R7452 AVDD.n2436 AVDD.n2372 21.9522
R7453 AVDD.n2380 AVDD.n2379 21.9522
R7454 AVDD.n2379 AVDD.n2377 21.9522
R7455 AVDD.n2413 AVDD.n2412 21.9522
R7456 AVDD.n2414 AVDD.n2413 21.9522
R7457 AVDD.n2395 AVDD.n2394 21.9522
R7458 AVDD.n2396 AVDD.n2395 21.9522
R7459 AVDD.n704 AVDD.n703 21.9522
R7460 AVDD.n703 AVDD.n702 21.9522
R7461 AVDD.n704 AVDD.n694 21.9522
R7462 AVDD.n702 AVDD.n694 21.9522
R7463 AVDD.n704 AVDD.n701 21.9522
R7464 AVDD.n702 AVDD.n701 21.9522
R7465 AVDD.n704 AVDD.n695 21.9522
R7466 AVDD.n702 AVDD.n695 21.9522
R7467 AVDD.n704 AVDD.n700 21.9522
R7468 AVDD.n702 AVDD.n700 21.9522
R7469 AVDD.n704 AVDD.n696 21.9522
R7470 AVDD.n702 AVDD.n696 21.9522
R7471 AVDD.n704 AVDD.n699 21.9522
R7472 AVDD.n702 AVDD.n699 21.9522
R7473 AVDD.n1073 AVDD.n1072 21.9522
R7474 AVDD.n1072 AVDD.n717 21.9522
R7475 AVDD.n1053 AVDD.n1052 21.9522
R7476 AVDD.n1054 AVDD.n1053 21.9522
R7477 AVDD.n1027 AVDD.n1026 21.9522
R7478 AVDD.n1028 AVDD.n1027 21.9522
R7479 AVDD.n971 AVDD.n970 21.9522
R7480 AVDD.n970 AVDD.n767 21.9522
R7481 AVDD.n1085 AVDD.n1084 21.9522
R7482 AVDD.n1086 AVDD.n1085 21.9522
R7483 AVDD.n1044 AVDD.n1043 21.9522
R7484 AVDD.n1045 AVDD.n1044 21.9522
R7485 AVDD.n1015 AVDD.n1014 21.9522
R7486 AVDD.n1014 AVDD.n1013 21.9522
R7487 AVDD.n2154 AVDD.n2153 21.9522
R7488 AVDD.n2155 AVDD.n2154 21.9522
R7489 AVDD.n2136 AVDD.n2135 21.9522
R7490 AVDD.n2137 AVDD.n2136 21.9522
R7491 AVDD.n2684 AVDD.n2120 21.9522
R7492 AVDD.n2685 AVDD.n2684 21.9522
R7493 AVDD.n2699 AVDD.n2698 21.9522
R7494 AVDD.n2698 AVDD.n2697 21.9522
R7495 AVDD.n2085 AVDD.n2084 21.9522
R7496 AVDD.n2086 AVDD.n2085 21.9522
R7497 AVDD.n2063 AVDD.n2062 21.9522
R7498 AVDD.n2064 AVDD.n2063 21.9522
R7499 AVDD.n2735 AVDD.n2047 21.9522
R7500 AVDD.n2736 AVDD.n2735 21.9522
R7501 AVDD.n2748 AVDD.n2033 21.9522
R7502 AVDD.n2749 AVDD.n2748 21.9522
R7503 AVDD.n2763 AVDD.n2762 21.9522
R7504 AVDD.n2762 AVDD.n2761 21.9522
R7505 AVDD.n2015 AVDD.n2003 21.9522
R7506 AVDD.n2016 AVDD.n2015 21.9522
R7507 AVDD.n2787 AVDD.n1989 21.9522
R7508 AVDD.n2788 AVDD.n2787 21.9522
R7509 AVDD.n2799 AVDD.n1969 21.9522
R7510 AVDD.n2800 AVDD.n2799 21.9522
R7511 AVDD.n2814 AVDD.n2813 21.9522
R7512 AVDD.n2813 AVDD.n2812 21.9522
R7513 AVDD.n1951 AVDD.n1939 21.9522
R7514 AVDD.n1952 AVDD.n1951 21.9522
R7515 AVDD.n3099 AVDD.n3098 21.8358
R7516 AVDD.n221 AVDD.n219 21.8358
R7517 AVDD.n3048 AVDD.n251 21.8358
R7518 AVDD.n3033 AVDD.n265 21.8358
R7519 AVDD.n2981 AVDD.n2980 21.8358
R7520 AVDD.n2951 AVDD.n339 21.8358
R7521 AVDD.n2936 AVDD.n359 21.8358
R7522 AVDD.n2906 AVDD.n2905 21.8358
R7523 AVDD.n416 AVDD.n414 21.8358
R7524 AVDD.n2855 AVDD.n444 21.8358
R7525 AVDD.n2840 AVDD.n457 21.8358
R7526 AVDD.n1350 AVDD.n1349 21.8358
R7527 AVDD.n1372 AVDD.n1371 21.8358
R7528 AVDD.n1680 AVDD.n1677 21.8358
R7529 AVDD.n1657 AVDD.n1656 21.8358
R7530 AVDD.n1604 AVDD.n1453 21.8358
R7531 AVDD.n1569 AVDD.n1566 21.8358
R7532 AVDD.n1547 AVDD.n1504 21.8358
R7533 AVDD.n2237 AVDD.n2235 21.8358
R7534 AVDD.n2263 AVDD.n2262 21.8358
R7535 AVDD.n2306 AVDD.n2305 21.8358
R7536 AVDD.n2326 AVDD.n2325 21.8358
R7537 AVDD.n1925 AVDD.n1924 21.8358
R7538 AVDD.n2391 AVDD.n2390 21.8358
R7539 AVDD.n2419 AVDD.n2418 21.8358
R7540 AVDD.n2456 AVDD.n2453 21.8358
R7541 AVDD.n2500 AVDD.n2499 21.8358
R7542 AVDD.n2548 AVDD.n2545 21.8358
R7543 AVDD.n2565 AVDD.n2564 21.8358
R7544 AVDD.n2614 AVDD.n2611 21.8358
R7545 AVDD.n2636 AVDD.n2635 21.8358
R7546 AVDD.n1880 AVDD.n519 21.8358
R7547 AVDD.n1865 AVDD.n533 21.8358
R7548 AVDD.n1833 AVDD.n1832 21.8358
R7549 AVDD.n1817 AVDD.n1164 21.8358
R7550 AVDD.n1786 AVDD.n1785 21.8358
R7551 AVDD.n1206 AVDD.n1204 21.8358
R7552 AVDD.n1920 AVDD.n505 21.8358
R7553 AVDD.n2823 AVDD.n1940 21.8358
R7554 AVDD.n1966 AVDD.n1958 21.8358
R7555 AVDD.n2772 AVDD.n2004 21.8358
R7556 AVDD.n2030 AVDD.n2022 21.8358
R7557 AVDD.n2720 AVDD.n2073 21.8358
R7558 AVDD.n2702 AVDD.n2099 21.8358
R7559 AVDD.n2669 AVDD.n2142 21.8358
R7560 AVDD.n2651 AVDD.n2168 21.8358
R7561 AVDD.n3286 AVDD.n3284 21.8358
R7562 AVDD.n3264 AVDD.n3263 21.8358
R7563 AVDD.n3229 AVDD.n3228 21.8358
R7564 AVDD.n3212 AVDD.n141 21.8358
R7565 AVDD.n3178 AVDD.n3177 21.8358
R7566 AVDD.n3158 AVDD.n168 21.8358
R7567 AVDD.n941 AVDD.n790 21.8358
R7568 AVDD.n920 AVDD.n919 21.8358
R7569 AVDD.n883 AVDD.n825 21.8358
R7570 AVDD.n864 AVDD.n840 21.8358
R7571 AVDD.n606 AVDD.n567 21.8358
R7572 AVDD.n623 AVDD.n584 21.8358
R7573 AVDD.n651 AVDD.n574 21.8358
R7574 AVDD.n668 AVDD.n588 21.8358
R7575 AVDD.n1096 AVDD.n718 21.4593
R7576 AVDD.n728 AVDD.n727 21.4593
R7577 AVDD.n1020 AVDD.t1 21.4192
R7578 AVDD.n1032 AVDD.n1031 20.7064
R7579 AVDD.n750 AVDD.n748 20.7064
R7580 AVDD.n202 AVDD.n199 20.3299
R7581 AVDD.n3079 AVDD.n223 20.3299
R7582 AVDD.n3049 AVDD.n246 20.3299
R7583 AVDD.n273 AVDD.n272 20.3299
R7584 AVDD.n296 AVDD.n293 20.3299
R7585 AVDD.n2976 AVDD.n316 20.3299
R7586 AVDD.n2952 AVDD.n336 20.3299
R7587 AVDD.n2932 AVDD.n2931 20.3299
R7588 AVDD.n401 AVDD.n399 20.3299
R7589 AVDD.n2882 AVDD.n418 20.3299
R7590 AVDD.n2856 AVDD.n442 20.3299
R7591 AVDD.n496 AVDD.n492 20.3299
R7592 AVDD.n1346 AVDD.n1332 20.3299
R7593 AVDD.n1375 AVDD.n1327 20.3299
R7594 AVDD.n1681 AVDD.n1394 20.3299
R7595 AVDD.n1653 AVDD.n1401 20.3299
R7596 AVDD.n1619 AVDD.n1444 20.3299
R7597 AVDD.n1601 AVDD.n1600 20.3299
R7598 AVDD.n1570 AVDD.n1492 20.3299
R7599 AVDD.n1543 AVDD.n1542 20.3299
R7600 AVDD.n3300 AVDD.n10 20.3299
R7601 AVDD.n2266 AVDD.n2229 20.3299
R7602 AVDD.n2302 AVDD.n2221 20.3299
R7603 AVDD.n2323 AVDD.n2322 20.3299
R7604 AVDD.n499 AVDD.n484 20.3299
R7605 AVDD.n2392 AVDD.n2389 20.3299
R7606 AVDD.n2423 AVDD.n2422 20.3299
R7607 AVDD.n2518 AVDD.n2516 20.3299
R7608 AVDD.n2498 AVDD.n2471 20.3299
R7609 AVDD.n2544 AVDD.n2543 20.3299
R7610 AVDD.n2569 AVDD.n2566 20.3299
R7611 AVDD.n2610 AVDD.n2609 20.3299
R7612 AVDD.n2196 AVDD.n2189 20.3299
R7613 AVDD.n1881 AVDD.n514 20.3299
R7614 AVDD.n541 AVDD.n540 20.3299
R7615 AVDD.n1147 AVDD.n1145 20.3299
R7616 AVDD.n1814 AVDD.n1813 20.3299
R7617 AVDD.n1193 AVDD.n1191 20.3299
R7618 AVDD.n1766 AVDD.n1208 20.3299
R7619 AVDD.n1919 AVDD.n506 20.3299
R7620 AVDD.n2824 AVDD.n476 20.3299
R7621 AVDD.n2803 AVDD.n1967 20.3299
R7622 AVDD.n2773 AVDD.n2000 20.3299
R7623 AVDD.n2752 AVDD.n2031 20.3299
R7624 AVDD.n2721 AVDD.n2059 20.3299
R7625 AVDD.n2701 AVDD.n2100 20.3299
R7626 AVDD.n2670 AVDD.n2132 20.3299
R7627 AVDD.n2650 AVDD.n2169 20.3299
R7628 AVDD.n3287 AVDD.n107 20.3299
R7629 AVDD.n3260 AVDD.n112 20.3299
R7630 AVDD.n3232 AVDD.n128 20.3299
R7631 AVDD.n3209 AVDD.n3208 20.3299
R7632 AVDD.n3181 AVDD.n161 20.3299
R7633 AVDD.n3151 AVDD.n3150 20.3299
R7634 AVDD.n942 AVDD.n786 20.3299
R7635 AVDD.n915 AVDD.n804 20.3299
R7636 AVDD.n887 AVDD.n886 20.3299
R7637 AVDD.n861 AVDD.n860 20.3299
R7638 AVDD.n603 AVDD.n579 20.3299
R7639 AVDD.n626 AVDD.n561 20.3299
R7640 AVDD.n648 AVDD.n571 20.3299
R7641 AVDD.n671 AVDD.n557 20.3299
R7642 AVDD.n1097 AVDD.n716 19.9534
R7643 AVDD.n1091 AVDD.n722 19.9534
R7644 AVDD.n1030 AVDD.n752 19.2005
R7645 AVDD.n1007 AVDD.n759 19.2005
R7646 AVDD.n3104 AVDD.n197 18.824
R7647 AVDD.n3078 AVDD.n224 18.824
R7648 AVDD.n3057 AVDD.n3056 18.824
R7649 AVDD.n3027 AVDD.n3026 18.824
R7650 AVDD.n3003 AVDD.n291 18.824
R7651 AVDD.n2975 AVDD.n320 18.824
R7652 AVDD.n2956 AVDD.n2955 18.824
R7653 AVDD.n363 AVDD.n361 18.824
R7654 AVDD.n2911 AVDD.n397 18.824
R7655 AVDD.n2881 AVDD.n419 18.824
R7656 AVDD.n2860 AVDD.n2859 18.824
R7657 AVDD.n1345 AVDD.n1334 18.824
R7658 AVDD.n1380 AVDD.n1379 18.824
R7659 AVDD.n1691 AVDD.n1688 18.824
R7660 AVDD.n1652 AVDD.n1402 18.824
R7661 AVDD.n1625 AVDD.n1622 18.824
R7662 AVDD.n1597 AVDD.n1596 18.824
R7663 AVDD.n1574 AVDD.n1573 18.824
R7664 AVDD.n1539 AVDD.n1538 18.824
R7665 AVDD.n3301 AVDD.n9 18.824
R7666 AVDD.n2270 AVDD.n2267 18.824
R7667 AVDD.n2301 AVDD.n2222 18.824
R7668 AVDD.n1902 AVDD.n489 18.824
R7669 AVDD.n2832 AVDD.n468 18.824
R7670 AVDD.n2421 AVDD.n2376 18.824
R7671 AVDD.n2519 AVDD.n2452 18.824
R7672 AVDD.n2480 AVDD.n2478 18.824
R7673 AVDD.n2541 AVDD.n2360 18.824
R7674 AVDD.n2570 AVDD.n2348 18.824
R7675 AVDD.n2607 AVDD.n2341 18.824
R7676 AVDD.n2210 AVDD.n2209 18.824
R7677 AVDD.n1889 AVDD.n1888 18.824
R7678 AVDD.n1859 AVDD.n1858 18.824
R7679 AVDD.n1838 AVDD.n1143 18.824
R7680 AVDD.n1170 AVDD.n1168 18.824
R7681 AVDD.n1791 AVDD.n1189 18.824
R7682 AVDD.n1765 AVDD.n1209 18.824
R7683 AVDD.n1905 AVDD.n508 18.824
R7684 AVDD.n2828 AVDD.n2827 18.824
R7685 AVDD.n2802 AVDD.n1968 18.824
R7686 AVDD.n2778 AVDD.n2777 18.824
R7687 AVDD.n2751 AVDD.n2032 18.824
R7688 AVDD.n2726 AVDD.n2725 18.824
R7689 AVDD.n2106 AVDD.n2105 18.824
R7690 AVDD.n2675 AVDD.n2674 18.824
R7691 AVDD.n2205 AVDD.n2171 18.824
R7692 AVDD.n106 AVDD.n99 18.824
R7693 AVDD.n3259 AVDD.n113 18.824
R7694 AVDD.n3236 AVDD.n3233 18.824
R7695 AVDD.n3205 AVDD.n3204 18.824
R7696 AVDD.n3185 AVDD.n3182 18.824
R7697 AVDD.n3147 AVDD.n3146 18.824
R7698 AVDD.n948 AVDD.n947 18.824
R7699 AVDD.n914 AVDD.n806 18.824
R7700 AVDD.n891 AVDD.n822 18.824
R7701 AVDD.n856 AVDD.n843 18.824
R7702 AVDD.n601 AVDD.n566 18.824
R7703 AVDD.n628 AVDD.n585 18.824
R7704 AVDD.n646 AVDD.n575 18.824
R7705 AVDD.n673 AVDD.n589 18.824
R7706 AVDD.n1101 AVDD.n1100 18.4476
R7707 AVDD.n1090 AVDD.n723 18.4476
R7708 AVDD.n1126 AVDD.t149 18.124
R7709 AVDD.n1024 AVDD.n1023 17.6946
R7710 AVDD.n1018 AVDD.n1017 17.6946
R7711 AVDD.n3105 AVDD.n193 17.3181
R7712 AVDD.n233 AVDD.n232 17.3181
R7713 AVDD.n245 AVDD.n243 17.3181
R7714 AVDD.n3022 AVDD.n274 17.3181
R7715 AVDD.n3004 AVDD.n286 17.3181
R7716 AVDD.n2972 AVDD.n2971 17.3181
R7717 AVDD.n335 AVDD.n333 17.3181
R7718 AVDD.n2926 AVDD.n365 17.3181
R7719 AVDD.n2912 AVDD.n380 17.3181
R7720 AVDD.n2878 AVDD.n2877 17.3181
R7721 AVDD.n2864 AVDD.n438 17.3181
R7722 AVDD.n1335 AVDD.n192 17.3181
R7723 AVDD.n1376 AVDD.n1321 17.3181
R7724 AVDD.n1692 AVDD.n1392 17.3181
R7725 AVDD.n1649 AVDD.n1648 17.3181
R7726 AVDD.n1626 AVDD.n1438 17.3181
R7727 AVDD.n1593 AVDD.n1461 17.3181
R7728 AVDD.n1577 AVDD.n1491 17.3181
R7729 AVDD.n1535 AVDD.n1506 17.3181
R7730 AVDD.n1519 AVDD.n1517 17.3181
R7731 AVDD.n2271 AVDD.n2227 17.3181
R7732 AVDD.n2297 AVDD.n2296 17.3181
R7733 AVDD.n1899 AVDD.n485 17.3181
R7734 AVDD.n2833 AVDD.n467 17.3181
R7735 AVDD.n2431 AVDD.n2430 17.3181
R7736 AVDD.n2451 AVDD.n2450 17.3181
R7737 AVDD.n2492 AVDD.n2491 17.3181
R7738 AVDD.n2533 AVDD.n2532 17.3181
R7739 AVDD.n2583 AVDD.n2582 17.3181
R7740 AVDD.n2599 AVDD.n2598 17.3181
R7741 AVDD.n2200 AVDD.n2190 17.3181
R7742 AVDD.n1893 AVDD.n512 17.3181
R7743 AVDD.n1854 AVDD.n542 17.3181
R7744 AVDD.n1839 AVDD.n553 17.3181
R7745 AVDD.n1808 AVDD.n1172 17.3181
R7746 AVDD.n1792 AVDD.n1187 17.3181
R7747 AVDD.n1761 AVDD.n1760 17.3181
R7748 AVDD.n1232 AVDD.n1228 17.3181
R7749 AVDD.n1744 AVDD.n1230 17.3181
R7750 AVDD.n1907 AVDD.n1896 17.3181
R7751 AVDD.n1934 AVDD.n475 17.3181
R7752 AVDD.n2797 AVDD.n2796 17.3181
R7753 AVDD.n1999 AVDD.n1998 17.3181
R7754 AVDD.n2746 AVDD.n2745 17.3181
R7755 AVDD.n2058 AVDD.n2057 17.3181
R7756 AVDD.n2695 AVDD.n2694 17.3181
R7757 AVDD.n2131 AVDD.n2130 17.3181
R7758 AVDD.n2203 AVDD.n2177 17.3181
R7759 AVDD.n3294 AVDD.n3293 17.3181
R7760 AVDD.n3256 AVDD.n3255 17.3181
R7761 AVDD.n3237 AVDD.n126 17.3181
R7762 AVDD.n3201 AVDD.n145 17.3181
R7763 AVDD.n3186 AVDD.n159 17.3181
R7764 AVDD.n3143 AVDD.n171 17.3181
R7765 AVDD.n185 AVDD.n177 17.3181
R7766 AVDD.n3124 AVDD.n3123 17.3181
R7767 AVDD.n966 AVDD.n784 17.3181
R7768 AVDD.n911 AVDD.n910 17.3181
R7769 AVDD.n892 AVDD.n819 17.3181
R7770 AVDD.n855 AVDD.n847 17.3181
R7771 AVDD.n598 AVDD.n580 17.3181
R7772 AVDD.n631 AVDD.n560 17.3181
R7773 AVDD.n643 AVDD.n570 17.3181
R7774 AVDD.n590 AVDD.n556 17.3181
R7775 AVDD.n974 AVDD.n780 16.9417
R7776 AVDD.n1102 AVDD.n707 16.9417
R7777 AVDD.n981 AVDD.n980 16.9417
R7778 AVDD.n1109 AVDD.n710 16.9417
R7779 AVDD.n1061 AVDD.t0 16.8059
R7780 AVDD.n766 AVDD.n754 16.1887
R7781 AVDD.n1132 AVDD.n683 16.1887
R7782 AVDD.n1002 AVDD.n758 16.1887
R7783 AVDD.n1129 AVDD.n1128 16.1887
R7784 AVDD.n3072 AVDD.n3071 15.8123
R7785 AVDD.n3062 AVDD.n241 15.8123
R7786 AVDD.n3021 AVDD.n278 15.8123
R7787 AVDD.n3012 AVDD.n3011 15.8123
R7788 AVDD.n324 AVDD.n322 15.8123
R7789 AVDD.n2961 AVDD.n331 15.8123
R7790 AVDD.n2925 AVDD.n366 15.8123
R7791 AVDD.n2916 AVDD.n2915 15.8123
R7792 AVDD.n425 AVDD.n423 15.8123
R7793 AVDD.n2865 AVDD.n437 15.8123
R7794 AVDD.n1387 AVDD.n1386 15.8123
R7795 AVDD.n1696 AVDD.n1695 15.8123
R7796 AVDD.n1645 AVDD.n1435 15.8123
R7797 AVDD.n1634 AVDD.n1633 15.8123
R7798 AVDD.n1592 AVDD.n1462 15.8123
R7799 AVDD.n1581 AVDD.n1578 15.8123
R7800 AVDD.n1534 AVDD.n1507 15.8123
R7801 AVDD.n1523 AVDD.n1522 15.8123
R7802 AVDD.n2277 AVDD.n2274 15.8123
R7803 AVDD.n2293 AVDD.n2292 15.8123
R7804 AVDD.n1901 AVDD.n488 15.8123
R7805 AVDD.n1929 AVDD.n1928 15.8123
R7806 AVDD.n2433 AVDD.n2432 15.8123
R7807 AVDD.n2449 AVDD.n2371 15.8123
R7808 AVDD.n2490 AVDD.n2481 15.8123
R7809 AVDD.n2534 AVDD.n2528 15.8123
R7810 AVDD.n2585 AVDD.n2584 15.8123
R7811 AVDD.n2600 AVDD.n2596 15.8123
R7812 AVDD.n2198 AVDD.n2195 15.8123
R7813 AVDD.n2639 AVDD.n2638 15.8123
R7814 AVDD.n1853 AVDD.n546 15.8123
R7815 AVDD.n1844 AVDD.n1843 15.8123
R7816 AVDD.n1807 AVDD.n1173 15.8123
R7817 AVDD.n1796 AVDD.n1795 15.8123
R7818 AVDD.n1220 AVDD.n1218 15.8123
R7819 AVDD.n1749 AVDD.n1226 15.8123
R7820 AVDD.n1743 AVDD.n1231 15.8123
R7821 AVDD.n1897 AVDD.n507 15.8123
R7822 AVDD.n1935 AVDD.n1933 15.8123
R7823 AVDD.n1984 AVDD.n1976 15.8123
R7824 AVDD.n2784 AVDD.n1991 15.8123
R7825 AVDD.n2042 AVDD.n2035 15.8123
R7826 AVDD.n2732 AVDD.n2049 15.8123
R7827 AVDD.n2115 AVDD.n2107 15.8123
R7828 AVDD.n2681 AVDD.n2122 15.8123
R7829 AVDD.n2178 AVDD.n2170 15.8123
R7830 AVDD.n2641 AVDD.n2176 15.8123
R7831 AVDD.n3252 AVDD.n3251 15.8123
R7832 AVDD.n3243 AVDD.n3240 15.8123
R7833 AVDD.n3200 AVDD.n146 15.8123
R7834 AVDD.n3190 AVDD.n3189 15.8123
R7835 AVDD.n3142 AVDD.n172 15.8123
R7836 AVDD.n3131 AVDD.n3130 15.8123
R7837 AVDD.n3120 AVDD.n3119 15.8123
R7838 AVDD.n956 AVDD.n955 15.8123
R7839 AVDD.n967 AVDD.n783 15.8123
R7840 AVDD.n906 AVDD.n808 15.8123
R7841 AVDD.n896 AVDD.n895 15.8123
R7842 AVDD.n850 AVDD.n774 15.8123
R7843 AVDD.n680 AVDD.n582 15.8123
R7844 AVDD.n596 AVDD.n565 15.8123
R7845 AVDD.n633 AVDD.n586 15.8123
R7846 AVDD.n641 AVDD.n576 15.8123
R7847 AVDD.n1140 AVDD.n1139 15.8123
R7848 AVDD.n986 AVDD.t130 15.4878
R7849 AVDD.n988 AVDD.n768 15.4358
R7850 AVDD.n1114 AVDD.n705 15.4358
R7851 AVDD.n984 AVDD.n771 15.4358
R7852 AVDD.n1108 AVDD.n711 15.4358
R7853 AVDD.n997 AVDD.n996 14.6829
R7854 AVDD.n697 AVDD.n688 14.6829
R7855 AVDD.n1003 AVDD.n1001 14.6829
R7856 AVDD.n692 AVDD.n685 14.6829
R7857 AVDD.n3067 AVDD.n234 14.3064
R7858 AVDD.n3063 AVDD.n238 14.3064
R7859 AVDD.n3018 AVDD.n3017 14.3064
R7860 AVDD.n285 AVDD.n283 14.3064
R7861 AVDD.n2966 AVDD.n326 14.3064
R7862 AVDD.n2962 AVDD.n327 14.3064
R7863 AVDD.n2922 AVDD.n2921 14.3064
R7864 AVDD.n379 AVDD.n377 14.3064
R7865 AVDD.n2872 AVDD.n427 14.3064
R7866 AVDD.n436 AVDD.n428 14.3064
R7867 AVDD.n1390 AVDD.n1320 14.3064
R7868 AVDD.n1699 AVDD.n1391 14.3064
R7869 AVDD.n1642 AVDD.n1641 14.3064
R7870 AVDD.n1637 AVDD.n1437 14.3064
R7871 AVDD.n1589 AVDD.n1588 14.3064
R7872 AVDD.n1582 AVDD.n1489 14.3064
R7873 AVDD.n1531 AVDD.n1530 14.3064
R7874 AVDD.n1526 AVDD.n1516 14.3064
R7875 AVDD.n2278 AVDD.n2225 14.3064
R7876 AVDD.n2289 AVDD.n2224 14.3064
R7877 AVDD.n1912 AVDD.n486 14.3064
R7878 AVDD.n1927 AVDD.n482 14.3064
R7879 AVDD.n2434 AVDD.n2373 14.3064
R7880 AVDD.n2442 AVDD.n2441 14.3064
R7881 AVDD.n2487 AVDD.n2486 14.3064
R7882 AVDD.n2527 AVDD.n2366 14.3064
R7883 AVDD.n2586 AVDD.n2346 14.3064
R7884 AVDD.n2595 AVDD.n2594 14.3064
R7885 AVDD.n2192 AVDD.n2191 14.3064
R7886 AVDD.n2193 AVDD.n2186 14.3064
R7887 AVDD.n1850 AVDD.n1849 14.3064
R7888 AVDD.n552 AVDD.n550 14.3064
R7889 AVDD.n1182 AVDD.n1181 14.3064
R7890 AVDD.n1800 AVDD.n1183 14.3064
R7891 AVDD.n1755 AVDD.n1222 14.3064
R7892 AVDD.n1750 AVDD.n1223 14.3064
R7893 AVDD.n1740 AVDD.n1739 14.3064
R7894 AVDD.n1731 AVDD.n1730 14.3064
R7895 AVDD.n1917 AVDD.n1916 14.3064
R7896 AVDD.n509 AVDD.n478 14.3064
R7897 AVDD.n2791 AVDD.n1985 14.3064
R7898 AVDD.n2785 AVDD.n1986 14.3064
R7899 AVDD.n2739 AVDD.n2043 14.3064
R7900 AVDD.n2733 AVDD.n2044 14.3064
R7901 AVDD.n2688 AVDD.n2116 14.3064
R7902 AVDD.n2682 AVDD.n2117 14.3064
R7903 AVDD.n2648 AVDD.n2647 14.3064
R7904 AVDD.n2180 AVDD.n2172 14.3064
R7905 AVDD.n3248 AVDD.n122 14.3064
R7906 AVDD.n3244 AVDD.n123 14.3064
R7907 AVDD.n157 AVDD.n154 14.3064
R7908 AVDD.n3193 AVDD.n158 14.3064
R7909 AVDD.n3139 AVDD.n3138 14.3064
R7910 AVDD.n3134 AVDD.n176 14.3064
R7911 AVDD.n3116 AVDD.n186 14.3064
R7912 AVDD.n3111 AVDD.n188 14.3064
R7913 AVDD.n959 AVDD.n953 14.3064
R7914 AVDD.n954 AVDD.n950 14.3064
R7915 AVDD.n905 AVDD.n811 14.3064
R7916 AVDD.n900 AVDD.n817 14.3064
R7917 AVDD.n678 AVDD.n563 14.3064
R7918 AVDD.n676 AVDD.n581 14.3064
R7919 AVDD.n636 AVDD.n559 14.3064
R7920 AVDD.n638 AVDD.n569 14.3064
R7921 AVDD.n990 AVDD.n989 13.9299
R7922 AVDD.n1116 AVDD.n1115 13.9299
R7923 AVDD.n983 AVDD.n772 13.9299
R7924 AVDD.n1120 AVDD.n691 13.9299
R7925 AVDD.n501 AVDD.n200 13.3358
R7926 AVDD.n989 AVDD.n765 13.177
R7927 AVDD.n1117 AVDD.n1116 13.177
R7928 AVDD.n772 AVDD.n761 13.177
R7929 AVDD.n1120 AVDD.n1119 13.177
R7930 AVDD.n3067 AVDD.n3066 12.8005
R7931 AVDD.n3066 AVDD.n238 12.8005
R7932 AVDD.n3017 AVDD.n281 12.8005
R7933 AVDD.n283 AVDD.n281 12.8005
R7934 AVDD.n2966 AVDD.n2965 12.8005
R7935 AVDD.n2965 AVDD.n327 12.8005
R7936 AVDD.n2921 AVDD.n375 12.8005
R7937 AVDD.n377 AVDD.n375 12.8005
R7938 AVDD.n2872 AVDD.n2871 12.8005
R7939 AVDD.n2871 AVDD.n428 12.8005
R7940 AVDD.n1700 AVDD.n1390 12.8005
R7941 AVDD.n1700 AVDD.n1699 12.8005
R7942 AVDD.n1641 AVDD.n1638 12.8005
R7943 AVDD.n1638 AVDD.n1637 12.8005
R7944 AVDD.n1588 AVDD.n1585 12.8005
R7945 AVDD.n1585 AVDD.n1489 12.8005
R7946 AVDD.n1530 AVDD.n1527 12.8005
R7947 AVDD.n1527 AVDD.n1526 12.8005
R7948 AVDD.n2288 AVDD.n2225 12.8005
R7949 AVDD.n2289 AVDD.n2288 12.8005
R7950 AVDD.n1912 AVDD.n487 12.8005
R7951 AVDD.n487 AVDD.n482 12.8005
R7952 AVDD.n2439 AVDD.n2373 12.8005
R7953 AVDD.n2441 AVDD.n2439 12.8005
R7954 AVDD.n2486 AVDD.n2485 12.8005
R7955 AVDD.n2485 AVDD.n2366 12.8005
R7956 AVDD.n2592 AVDD.n2346 12.8005
R7957 AVDD.n2594 AVDD.n2592 12.8005
R7958 AVDD.n2194 AVDD.n2192 12.8005
R7959 AVDD.n2194 AVDD.n2193 12.8005
R7960 AVDD.n1849 AVDD.n548 12.8005
R7961 AVDD.n550 AVDD.n548 12.8005
R7962 AVDD.n1801 AVDD.n1182 12.8005
R7963 AVDD.n1801 AVDD.n1800 12.8005
R7964 AVDD.n1755 AVDD.n1754 12.8005
R7965 AVDD.n1754 AVDD.n1223 12.8005
R7966 AVDD.n1739 AVDD.n1728 12.8005
R7967 AVDD.n1731 AVDD.n1728 12.8005
R7968 AVDD.n1916 AVDD.n510 12.8005
R7969 AVDD.n510 AVDD.n509 12.8005
R7970 AVDD.n2791 AVDD.n2790 12.8005
R7971 AVDD.n2790 AVDD.n1986 12.8005
R7972 AVDD.n2739 AVDD.n2738 12.8005
R7973 AVDD.n2738 AVDD.n2044 12.8005
R7974 AVDD.n2688 AVDD.n2687 12.8005
R7975 AVDD.n2687 AVDD.n2117 12.8005
R7976 AVDD.n2647 AVDD.n2174 12.8005
R7977 AVDD.n2180 AVDD.n2174 12.8005
R7978 AVDD.n3248 AVDD.n3247 12.8005
R7979 AVDD.n3247 AVDD.n123 12.8005
R7980 AVDD.n3194 AVDD.n157 12.8005
R7981 AVDD.n3194 AVDD.n3193 12.8005
R7982 AVDD.n3138 AVDD.n3135 12.8005
R7983 AVDD.n3135 AVDD.n3134 12.8005
R7984 AVDD.n3116 AVDD.n3115 12.8005
R7985 AVDD.n3115 AVDD.n188 12.8005
R7986 AVDD.n959 AVDD.n958 12.8005
R7987 AVDD.n958 AVDD.n950 12.8005
R7988 AVDD.n901 AVDD.n811 12.8005
R7989 AVDD.n901 AVDD.n900 12.8005
R7990 AVDD.n678 AVDD.n564 12.8005
R7991 AVDD.n676 AVDD.n564 12.8005
R7992 AVDD.n636 AVDD.n577 12.8005
R7993 AVDD.n638 AVDD.n577 12.8005
R7994 AVDD.n997 AVDD.n765 12.424
R7995 AVDD.n1117 AVDD.n688 12.424
R7996 AVDD.n1001 AVDD.n761 12.424
R7997 AVDD.n1119 AVDD.n692 12.424
R7998 AVDD.n1079 AVDD.t2 12.1927
R7999 AVDD.n990 AVDD.n988 11.6711
R8000 AVDD.n1115 AVDD.n1114 11.6711
R8001 AVDD.n984 AVDD.n983 11.6711
R8002 AVDD.n711 AVDD.n691 11.6711
R8003 AVDD.n3071 AVDD.n234 11.2946
R8004 AVDD.n3063 AVDD.n3062 11.2946
R8005 AVDD.n3018 AVDD.n278 11.2946
R8006 AVDD.n3012 AVDD.n285 11.2946
R8007 AVDD.n326 AVDD.n324 11.2946
R8008 AVDD.n2962 AVDD.n2961 11.2946
R8009 AVDD.n2922 AVDD.n366 11.2946
R8010 AVDD.n2916 AVDD.n379 11.2946
R8011 AVDD.n427 AVDD.n425 11.2946
R8012 AVDD.n437 AVDD.n436 11.2946
R8013 AVDD.n1387 AVDD.n1320 11.2946
R8014 AVDD.n1696 AVDD.n1391 11.2946
R8015 AVDD.n1642 AVDD.n1435 11.2946
R8016 AVDD.n1634 AVDD.n1437 11.2946
R8017 AVDD.n1589 AVDD.n1462 11.2946
R8018 AVDD.n1582 AVDD.n1581 11.2946
R8019 AVDD.n1531 AVDD.n1507 11.2946
R8020 AVDD.n1523 AVDD.n1516 11.2946
R8021 AVDD.n2278 AVDD.n2277 11.2946
R8022 AVDD.n2292 AVDD.n2224 11.2946
R8023 AVDD.n1901 AVDD.n486 11.2946
R8024 AVDD.n1929 AVDD.n1927 11.2946
R8025 AVDD.n2434 AVDD.n2433 11.2946
R8026 AVDD.n2442 AVDD.n2371 11.2946
R8027 AVDD.n2487 AVDD.n2481 11.2946
R8028 AVDD.n2528 AVDD.n2527 11.2946
R8029 AVDD.n2586 AVDD.n2585 11.2946
R8030 AVDD.n2596 AVDD.n2595 11.2946
R8031 AVDD.n2198 AVDD.n2191 11.2946
R8032 AVDD.n2639 AVDD.n2186 11.2946
R8033 AVDD.n1850 AVDD.n546 11.2946
R8034 AVDD.n1844 AVDD.n552 11.2946
R8035 AVDD.n1181 AVDD.n1173 11.2946
R8036 AVDD.n1796 AVDD.n1183 11.2946
R8037 AVDD.n1222 AVDD.n1220 11.2946
R8038 AVDD.n1750 AVDD.n1749 11.2946
R8039 AVDD.n1740 AVDD.n1231 11.2946
R8040 AVDD.n1730 AVDD.n194 11.2946
R8041 AVDD.n1917 AVDD.n1897 11.2946
R8042 AVDD.n1933 AVDD.n478 11.2946
R8043 AVDD.n1985 AVDD.n1984 11.2946
R8044 AVDD.n2785 AVDD.n2784 11.2946
R8045 AVDD.n2043 AVDD.n2042 11.2946
R8046 AVDD.n2733 AVDD.n2732 11.2946
R8047 AVDD.n2116 AVDD.n2115 11.2946
R8048 AVDD.n2682 AVDD.n2681 11.2946
R8049 AVDD.n2648 AVDD.n2178 11.2946
R8050 AVDD.n2641 AVDD.n2172 11.2946
R8051 AVDD.n3251 AVDD.n122 11.2946
R8052 AVDD.n3244 AVDD.n3243 11.2946
R8053 AVDD.n154 AVDD.n146 11.2946
R8054 AVDD.n3190 AVDD.n158 11.2946
R8055 AVDD.n3139 AVDD.n172 11.2946
R8056 AVDD.n3131 AVDD.n176 11.2946
R8057 AVDD.n3119 AVDD.n186 11.2946
R8058 AVDD.n3111 AVDD.n3110 11.2946
R8059 AVDD.n955 AVDD.n953 11.2946
R8060 AVDD.n954 AVDD.n783 11.2946
R8061 AVDD.n906 AVDD.n905 11.2946
R8062 AVDD.n896 AVDD.n817 11.2946
R8063 AVDD.n680 AVDD.n563 11.2946
R8064 AVDD.n596 AVDD.n581 11.2946
R8065 AVDD.n633 AVDD.n559 11.2946
R8066 AVDD.n641 AVDD.n569 11.2946
R8067 AVDD.n996 AVDD.n766 10.9181
R8068 AVDD.n697 AVDD.n683 10.9181
R8069 AVDD.n1003 AVDD.n1002 10.9181
R8070 AVDD.n1128 AVDD.n685 10.9181
R8071 AVDD.n1094 AVDD.t2 10.2156
R8072 AVDD.n2998 AVDD.n2997 10.1652
R8073 AVDD.n1618 AVDD.n298 10.1652
R8074 AVDD.n780 AVDD.n768 10.1652
R8075 AVDD.n707 AVDD.n705 10.1652
R8076 AVDD.n980 AVDD.n771 10.1652
R8077 AVDD.n1109 AVDD.n1108 10.1652
R8078 AVDD.n3297 AVDD.n13 9.89974
R8079 AVDD.n3072 AVDD.n233 9.78874
R8080 AVDD.n243 AVDD.n241 9.78874
R8081 AVDD.n3022 AVDD.n3021 9.78874
R8082 AVDD.n3011 AVDD.n286 9.78874
R8083 AVDD.n2971 AVDD.n322 9.78874
R8084 AVDD.n333 AVDD.n331 9.78874
R8085 AVDD.n2926 AVDD.n2925 9.78874
R8086 AVDD.n2915 AVDD.n380 9.78874
R8087 AVDD.n2877 AVDD.n423 9.78874
R8088 AVDD.n2865 AVDD.n2864 9.78874
R8089 AVDD.n1386 AVDD.n1321 9.78874
R8090 AVDD.n1695 AVDD.n1392 9.78874
R8091 AVDD.n1648 AVDD.n1645 9.78874
R8092 AVDD.n1633 AVDD.n1438 9.78874
R8093 AVDD.n1593 AVDD.n1592 9.78874
R8094 AVDD.n1578 AVDD.n1577 9.78874
R8095 AVDD.n1535 AVDD.n1534 9.78874
R8096 AVDD.n1522 AVDD.n1519 9.78874
R8097 AVDD.n2274 AVDD.n2227 9.78874
R8098 AVDD.n2296 AVDD.n2293 9.78874
R8099 AVDD.n1899 AVDD.n488 9.78874
R8100 AVDD.n1928 AVDD.n467 9.78874
R8101 AVDD.n2432 AVDD.n2431 9.78874
R8102 AVDD.n2450 AVDD.n2449 9.78874
R8103 AVDD.n2491 AVDD.n2490 9.78874
R8104 AVDD.n2534 AVDD.n2533 9.78874
R8105 AVDD.n2584 AVDD.n2583 9.78874
R8106 AVDD.n2600 AVDD.n2599 9.78874
R8107 AVDD.n2200 AVDD.n2195 9.78874
R8108 AVDD.n2638 AVDD.n2187 9.78874
R8109 AVDD.n1894 AVDD.n1893 9.78874
R8110 AVDD.n1854 AVDD.n1853 9.78874
R8111 AVDD.n1843 AVDD.n553 9.78874
R8112 AVDD.n1808 AVDD.n1807 9.78874
R8113 AVDD.n1795 AVDD.n1187 9.78874
R8114 AVDD.n1760 AVDD.n1218 9.78874
R8115 AVDD.n1228 AVDD.n1226 9.78874
R8116 AVDD.n1744 AVDD.n1743 9.78874
R8117 AVDD.n1907 AVDD.n507 9.78874
R8118 AVDD.n1935 AVDD.n1934 9.78874
R8119 AVDD.n2796 AVDD.n1976 9.78874
R8120 AVDD.n1998 AVDD.n1991 9.78874
R8121 AVDD.n2745 AVDD.n2035 9.78874
R8122 AVDD.n2057 AVDD.n2049 9.78874
R8123 AVDD.n2694 AVDD.n2107 9.78874
R8124 AVDD.n2130 AVDD.n2122 9.78874
R8125 AVDD.n2203 AVDD.n2170 9.78874
R8126 AVDD.n2176 AVDD.n2175 9.78874
R8127 AVDD.n3294 AVDD.n98 9.78874
R8128 AVDD.n3255 AVDD.n3252 9.78874
R8129 AVDD.n3240 AVDD.n126 9.78874
R8130 AVDD.n3201 AVDD.n3200 9.78874
R8131 AVDD.n3189 AVDD.n159 9.78874
R8132 AVDD.n3143 AVDD.n3142 9.78874
R8133 AVDD.n3130 AVDD.n177 9.78874
R8134 AVDD.n3123 AVDD.n3120 9.78874
R8135 AVDD.n956 AVDD.n779 9.78874
R8136 AVDD.n967 AVDD.n966 9.78874
R8137 AVDD.n910 AVDD.n808 9.78874
R8138 AVDD.n895 AVDD.n819 9.78874
R8139 AVDD.n850 AVDD.n847 9.78874
R8140 AVDD.n1134 AVDD.n582 9.78874
R8141 AVDD.n598 AVDD.n565 9.78874
R8142 AVDD.n631 AVDD.n586 9.78874
R8143 AVDD.n643 AVDD.n576 9.78874
R8144 AVDD.n1140 AVDD.n590 9.78874
R8145 AVDD.n1023 AVDD.n754 9.41227
R8146 AVDD.n1133 AVDD.n1132 9.41227
R8147 AVDD.n1018 AVDD.n758 9.41227
R8148 AVDD.n1129 AVDD.n591 9.41227
R8149 AVDD.n1936 AVDD.n1935 9.3005
R8150 AVDD.n1937 AVDD.n475 9.3005
R8151 AVDD.n2827 AVDD.n2826 9.3005
R8152 AVDD.n2825 AVDD.n2824 9.3005
R8153 AVDD.n1950 AVDD.n1940 9.3005
R8154 AVDD.n1953 AVDD.n1948 9.3005
R8155 AVDD.n2816 AVDD.n2815 9.3005
R8156 AVDD.n2790 AVDD.n2789 9.3005
R8157 AVDD.n2786 AVDD.n2785 9.3005
R8158 AVDD.n2001 AVDD.n1991 9.3005
R8159 AVDD.n2002 AVDD.n1999 9.3005
R8160 AVDD.n2777 AVDD.n2776 9.3005
R8161 AVDD.n2774 AVDD.n2773 9.3005
R8162 AVDD.n2014 AVDD.n2004 9.3005
R8163 AVDD.n2017 AVDD.n2012 9.3005
R8164 AVDD.n2765 AVDD.n2764 9.3005
R8165 AVDD.n2738 AVDD.n2737 9.3005
R8166 AVDD.n2734 AVDD.n2733 9.3005
R8167 AVDD.n2061 AVDD.n2049 9.3005
R8168 AVDD.n2060 AVDD.n2058 9.3005
R8169 AVDD.n2725 AVDD.n2724 9.3005
R8170 AVDD.n2722 AVDD.n2721 9.3005
R8171 AVDD.n2073 AVDD.n2072 9.3005
R8172 AVDD.n2083 AVDD.n2081 9.3005
R8173 AVDD.n2713 AVDD.n2712 9.3005
R8174 AVDD.n2687 AVDD.n2686 9.3005
R8175 AVDD.n2683 AVDD.n2682 9.3005
R8176 AVDD.n2134 AVDD.n2122 9.3005
R8177 AVDD.n2133 AVDD.n2131 9.3005
R8178 AVDD.n2674 AVDD.n2673 9.3005
R8179 AVDD.n2671 AVDD.n2670 9.3005
R8180 AVDD.n2142 AVDD.n2141 9.3005
R8181 AVDD.n2152 AVDD.n2150 9.3005
R8182 AVDD.n2662 AVDD.n2661 9.3005
R8183 AVDD.n2403 AVDD.n1955 9.3005
R8184 AVDD.n2811 AVDD.n2810 9.3005
R8185 AVDD.n1958 AVDD.n1956 9.3005
R8186 AVDD.n1971 AVDD.n1967 9.3005
R8187 AVDD.n2802 AVDD.n2801 9.3005
R8188 AVDD.n2798 AVDD.n2797 9.3005
R8189 AVDD.n1987 AVDD.n1976 9.3005
R8190 AVDD.n1988 AVDD.n1985 9.3005
R8191 AVDD.n2464 AVDD.n2019 9.3005
R8192 AVDD.n2760 AVDD.n2759 9.3005
R8193 AVDD.n2022 AVDD.n2020 9.3005
R8194 AVDD.n2066 AVDD.n2031 9.3005
R8195 AVDD.n2751 AVDD.n2750 9.3005
R8196 AVDD.n2747 AVDD.n2746 9.3005
R8197 AVDD.n2045 AVDD.n2035 9.3005
R8198 AVDD.n2046 AVDD.n2043 9.3005
R8199 AVDD.n2710 AVDD.n2709 9.3005
R8200 AVDD.n2089 AVDD.n2087 9.3005
R8201 AVDD.n2101 AVDD.n2099 9.3005
R8202 AVDD.n2701 AVDD.n2700 9.3005
R8203 AVDD.n2105 AVDD.n2103 9.3005
R8204 AVDD.n2696 AVDD.n2695 9.3005
R8205 AVDD.n2118 AVDD.n2107 9.3005
R8206 AVDD.n2119 AVDD.n2116 9.3005
R8207 AVDD.n2659 AVDD.n2658 9.3005
R8208 AVDD.n2158 AVDD.n2156 9.3005
R8209 AVDD.n2637 AVDD.n2194 9.3005
R8210 AVDD.n2637 AVDD.n2186 9.3005
R8211 AVDD.n2638 AVDD.n2637 9.3005
R8212 AVDD.n2313 AVDD.n2312 9.3005
R8213 AVDD.n2311 AVDD.n2310 9.3005
R8214 AVDD.n2306 AVDD.n2220 9.3005
R8215 AVDD.n2299 AVDD.n2221 9.3005
R8216 AVDD.n2301 AVDD.n2300 9.3005
R8217 AVDD.n2298 AVDD.n2297 9.3005
R8218 AVDD.n2293 AVDD.n2223 9.3005
R8219 AVDD.n2281 AVDD.n2224 9.3005
R8220 AVDD.n2288 AVDD.n2287 9.3005
R8221 AVDD.n2246 AVDD.n2245 9.3005
R8222 AVDD.n2234 AVDD.n2233 9.3005
R8223 AVDD.n2237 AVDD.n2236 9.3005
R8224 AVDD.n10 AVDD.n8 9.3005
R8225 AVDD.n3302 AVDD.n3301 9.3005
R8226 AVDD.n1517 AVDD.n7 9.3005
R8227 AVDD.n1522 AVDD.n1521 9.3005
R8228 AVDD.n1520 AVDD.n1516 9.3005
R8229 AVDD.n1527 AVDD.n1515 9.3005
R8230 AVDD.n1555 AVDD.n1554 9.3005
R8231 AVDD.n1560 AVDD.n1559 9.3005
R8232 AVDD.n1566 AVDD.n1565 9.3005
R8233 AVDD.n1571 AVDD.n1570 9.3005
R8234 AVDD.n1573 AVDD.n1572 9.3005
R8235 AVDD.n1493 AVDD.n1491 9.3005
R8236 AVDD.n1578 AVDD.n1490 9.3005
R8237 AVDD.n1583 AVDD.n1582 9.3005
R8238 AVDD.n1585 AVDD.n1584 9.3005
R8239 AVDD.n1612 AVDD.n1611 9.3005
R8240 AVDD.n1616 AVDD.n1615 9.3005
R8241 AVDD.n1617 AVDD.n298 9.3005
R8242 AVDD.n1620 AVDD.n1619 9.3005
R8243 AVDD.n1622 AVDD.n1621 9.3005
R8244 AVDD.n1627 AVDD.n1626 9.3005
R8245 AVDD.n1633 AVDD.n1632 9.3005
R8246 AVDD.n1439 AVDD.n1437 9.3005
R8247 AVDD.n1638 AVDD.n1436 9.3005
R8248 AVDD.n1670 AVDD.n1398 9.3005
R8249 AVDD.n1675 AVDD.n1674 9.3005
R8250 AVDD.n1677 AVDD.n1676 9.3005
R8251 AVDD.n1682 AVDD.n1681 9.3005
R8252 AVDD.n1688 AVDD.n1687 9.3005
R8253 AVDD.n1693 AVDD.n1692 9.3005
R8254 AVDD.n1695 AVDD.n1694 9.3005
R8255 AVDD.n1391 AVDD.n1319 9.3005
R8256 AVDD.n1701 AVDD.n1700 9.3005
R8257 AVDD.n1358 AVDD.n1357 9.3005
R8258 AVDD.n1355 AVDD.n1354 9.3005
R8259 AVDD.n1350 AVDD.n1331 9.3005
R8260 AVDD.n1338 AVDD.n1332 9.3005
R8261 AVDD.n1345 AVDD.n1344 9.3005
R8262 AVDD.n1336 AVDD.n1335 9.3005
R8263 AVDD.n2649 AVDD.n2174 9.3005
R8264 AVDD.n2649 AVDD.n2172 9.3005
R8265 AVDD.n2649 AVDD.n2176 9.3005
R8266 AVDD.n1363 AVDD.n1329 9.3005
R8267 AVDD.n1368 AVDD.n1367 9.3005
R8268 AVDD.n1371 AVDD.n1370 9.3005
R8269 AVDD.n1327 AVDD.n1326 9.3005
R8270 AVDD.n1381 AVDD.n1380 9.3005
R8271 AVDD.n1376 AVDD.n1322 9.3005
R8272 AVDD.n1386 AVDD.n1385 9.3005
R8273 AVDD.n1320 AVDD.n1318 9.3005
R8274 AVDD.n1665 AVDD.n1664 9.3005
R8275 AVDD.n1662 AVDD.n1661 9.3005
R8276 AVDD.n1657 AVDD.n1400 9.3005
R8277 AVDD.n1403 AVDD.n1401 9.3005
R8278 AVDD.n1652 AVDD.n1651 9.3005
R8279 AVDD.n1650 AVDD.n1649 9.3005
R8280 AVDD.n1645 AVDD.n1644 9.3005
R8281 AVDD.n1643 AVDD.n1642 9.3005
R8282 AVDD.n1610 AVDD.n1609 9.3005
R8283 AVDD.n1454 AVDD.n1452 9.3005
R8284 AVDD.n1604 AVDD.n1603 9.3005
R8285 AVDD.n1602 AVDD.n1601 9.3005
R8286 AVDD.n1597 AVDD.n1460 9.3005
R8287 AVDD.n1463 AVDD.n1461 9.3005
R8288 AVDD.n1592 AVDD.n1591 9.3005
R8289 AVDD.n1590 AVDD.n1589 9.3005
R8290 AVDD.n1553 AVDD.n1552 9.3005
R8291 AVDD.n1503 AVDD.n1499 9.3005
R8292 AVDD.n1547 AVDD.n1546 9.3005
R8293 AVDD.n1544 AVDD.n1543 9.3005
R8294 AVDD.n1539 AVDD.n1505 9.3005
R8295 AVDD.n1508 AVDD.n1506 9.3005
R8296 AVDD.n1534 AVDD.n1533 9.3005
R8297 AVDD.n1532 AVDD.n1531 9.3005
R8298 AVDD.n2253 AVDD.n2252 9.3005
R8299 AVDD.n2258 AVDD.n2257 9.3005
R8300 AVDD.n2262 AVDD.n2261 9.3005
R8301 AVDD.n2259 AVDD.n2229 9.3005
R8302 AVDD.n2267 AVDD.n2228 9.3005
R8303 AVDD.n2272 AVDD.n2271 9.3005
R8304 AVDD.n2274 AVDD.n2273 9.3005
R8305 AVDD.n2279 AVDD.n2278 9.3005
R8306 AVDD.n2318 AVDD.n2218 9.3005
R8307 AVDD.n2331 AVDD.n2330 9.3005
R8308 AVDD.n2326 AVDD.n2213 9.3005
R8309 AVDD.n2323 AVDD.n2215 9.3005
R8310 AVDD.n2321 AVDD.n2320 9.3005
R8311 AVDD.n2637 AVDD.n2191 9.3005
R8312 AVDD.n2637 AVDD.n2195 9.3005
R8313 AVDD.n2637 AVDD.n2190 9.3005
R8314 AVDD.n2637 AVDD.n2210 9.3005
R8315 AVDD.n2637 AVDD.n2189 9.3005
R8316 AVDD.n2637 AVDD.n2636 9.3005
R8317 AVDD.n2649 AVDD.n2168 9.3005
R8318 AVDD.n2650 AVDD.n2649 9.3005
R8319 AVDD.n2649 AVDD.n2171 9.3005
R8320 AVDD.n2649 AVDD.n2177 9.3005
R8321 AVDD.n2649 AVDD.n2170 9.3005
R8322 AVDD.n2649 AVDD.n2648 9.3005
R8323 AVDD.n3109 AVDD.n191 9.3005
R8324 AVDD.n3112 AVDD.n3111 9.3005
R8325 AVDD.n3115 AVDD.n3114 9.3005
R8326 AVDD.n3125 AVDD.n3124 9.3005
R8327 AVDD.n185 AVDD.n181 9.3005
R8328 AVDD.n3130 AVDD.n3129 9.3005
R8329 AVDD.n179 AVDD.n176 9.3005
R8330 AVDD.n3135 AVDD.n175 9.3005
R8331 AVDD.n3170 AVDD.n165 9.3005
R8332 AVDD.n3175 AVDD.n3174 9.3005
R8333 AVDD.n3177 AVDD.n3176 9.3005
R8334 AVDD.n163 AVDD.n161 9.3005
R8335 AVDD.n3182 AVDD.n160 9.3005
R8336 AVDD.n3187 AVDD.n3186 9.3005
R8337 AVDD.n3189 AVDD.n3188 9.3005
R8338 AVDD.n158 AVDD.n153 9.3005
R8339 AVDD.n3195 AVDD.n3194 9.3005
R8340 AVDD.n3223 AVDD.n3222 9.3005
R8341 AVDD.n136 AVDD.n132 9.3005
R8342 AVDD.n3228 AVDD.n3227 9.3005
R8343 AVDD.n130 AVDD.n128 9.3005
R8344 AVDD.n3233 AVDD.n127 9.3005
R8345 AVDD.n3238 AVDD.n3237 9.3005
R8346 AVDD.n3240 AVDD.n3239 9.3005
R8347 AVDD.n3245 AVDD.n3244 9.3005
R8348 AVDD.n3247 AVDD.n3246 9.3005
R8349 AVDD.n3277 AVDD.n109 9.3005
R8350 AVDD.n3282 AVDD.n3281 9.3005
R8351 AVDD.n3284 AVDD.n3283 9.3005
R8352 AVDD.n3288 AVDD.n3287 9.3005
R8353 AVDD.n106 AVDD.n102 9.3005
R8354 AVDD.n3293 AVDD.n3292 9.3005
R8355 AVDD.n2173 AVDD.n98 9.3005
R8356 AVDD.n3272 AVDD.n3271 9.3005
R8357 AVDD.n3269 AVDD.n3268 9.3005
R8358 AVDD.n3264 AVDD.n111 9.3005
R8359 AVDD.n114 AVDD.n112 9.3005
R8360 AVDD.n3259 AVDD.n3258 9.3005
R8361 AVDD.n3257 AVDD.n3256 9.3005
R8362 AVDD.n3252 AVDD.n121 9.3005
R8363 AVDD.n124 AVDD.n122 9.3005
R8364 AVDD.n3217 AVDD.n135 9.3005
R8365 AVDD.n143 AVDD.n140 9.3005
R8366 AVDD.n3212 AVDD.n3211 9.3005
R8367 AVDD.n3210 AVDD.n3209 9.3005
R8368 AVDD.n3205 AVDD.n144 9.3005
R8369 AVDD.n148 AVDD.n145 9.3005
R8370 AVDD.n3200 AVDD.n3199 9.3005
R8371 AVDD.n154 AVDD.n150 9.3005
R8372 AVDD.n3165 AVDD.n3164 9.3005
R8373 AVDD.n3163 AVDD.n3162 9.3005
R8374 AVDD.n3158 AVDD.n3157 9.3005
R8375 AVDD.n3152 AVDD.n3151 9.3005
R8376 AVDD.n3147 AVDD.n170 9.3005
R8377 AVDD.n174 AVDD.n171 9.3005
R8378 AVDD.n3142 AVDD.n3141 9.3005
R8379 AVDD.n3140 AVDD.n3139 9.3005
R8380 AVDD.n3120 AVDD.n184 9.3005
R8381 AVDD.n189 AVDD.n186 9.3005
R8382 AVDD.n1004 AVDD.n1003 9.3005
R8383 AVDD.n1005 AVDD.n758 9.3005
R8384 AVDD.n1017 AVDD.n1016 9.3005
R8385 AVDD.n1008 AVDD.n1007 9.3005
R8386 AVDD.n1012 AVDD.n748 9.3005
R8387 AVDD.n1038 AVDD.n747 9.3005
R8388 AVDD.n1042 AVDD.n1041 9.3005
R8389 AVDD.n746 AVDD.n745 9.3005
R8390 AVDD.n1108 AVDD.n1107 9.3005
R8391 AVDD.n712 AVDD.n710 9.3005
R8392 AVDD.n1090 AVDD.n1089 9.3005
R8393 AVDD.n1087 AVDD.n722 9.3005
R8394 AVDD.n728 AVDD.n724 9.3005
R8395 AVDD.n1083 AVDD.n1082 9.3005
R8396 AVDD.n1047 AVDD.n1046 9.3005
R8397 AVDD.n982 AVDD.n761 9.3005
R8398 AVDD.n877 AVDD.n876 9.3005
R8399 AVDD.n831 AVDD.n830 9.3005
R8400 AVDD.n884 AVDD.n883 9.3005
R8401 AVDD.n886 AVDD.n885 9.3005
R8402 AVDD.n826 AVDD.n822 9.3005
R8403 AVDD.n893 AVDD.n892 9.3005
R8404 AVDD.n895 AVDD.n894 9.3005
R8405 AVDD.n817 AVDD.n816 9.3005
R8406 AVDD.n902 AVDD.n901 9.3005
R8407 AVDD.n934 AVDD.n933 9.3005
R8408 AVDD.n936 AVDD.n935 9.3005
R8409 AVDD.n790 AVDD.n789 9.3005
R8410 AVDD.n943 AVDD.n942 9.3005
R8411 AVDD.n947 AVDD.n946 9.3005
R8412 AVDD.n784 AVDD.n782 9.3005
R8413 AVDD.n968 AVDD.n967 9.3005
R8414 AVDD.n983 AVDD.n982 9.3005
R8415 AVDD.n982 AVDD.n771 9.3005
R8416 AVDD.n982 AVDD.n981 9.3005
R8417 AVDD.n851 AVDD.n850 9.3005
R8418 AVDD.n855 AVDD.n854 9.3005
R8419 AVDD.n848 AVDD.n843 9.3005
R8420 AVDD.n862 AVDD.n861 9.3005
R8421 AVDD.n864 AVDD.n863 9.3005
R8422 AVDD.n838 AVDD.n836 9.3005
R8423 AVDD.n873 AVDD.n872 9.3005
R8424 AVDD.n905 AVDD.n904 9.3005
R8425 AVDD.n812 AVDD.n808 9.3005
R8426 AVDD.n912 AVDD.n911 9.3005
R8427 AVDD.n914 AVDD.n913 9.3005
R8428 AVDD.n804 AVDD.n803 9.3005
R8429 AVDD.n921 AVDD.n920 9.3005
R8430 AVDD.n925 AVDD.n924 9.3005
R8431 AVDD.n800 AVDD.n798 9.3005
R8432 AVDD.n957 AVDD.n954 9.3005
R8433 AVDD.n958 AVDD.n957 9.3005
R8434 AVDD.n993 AVDD.n765 9.3005
R8435 AVDD.n996 AVDD.n995 9.3005
R8436 AVDD.n994 AVDD.n754 9.3005
R8437 AVDD.n1025 AVDD.n1024 9.3005
R8438 AVDD.n1030 AVDD.n1029 9.3005
R8439 AVDD.n1031 AVDD.n735 9.3005
R8440 AVDD.n1066 AVDD.n1065 9.3005
R8441 AVDD.n738 AVDD.n736 9.3005
R8442 AVDD.n1056 AVDD.n1055 9.3005
R8443 AVDD.n957 AVDD.n953 9.3005
R8444 AVDD.n957 AVDD.n956 9.3005
R8445 AVDD.n974 AVDD.n973 9.3005
R8446 AVDD.n969 AVDD.n768 9.3005
R8447 AVDD.n991 AVDD.n990 9.3005
R8448 AVDD.n734 AVDD.n732 9.3005
R8449 AVDD.n1075 AVDD.n1074 9.3005
R8450 AVDD.n1071 AVDD.n718 9.3005
R8451 AVDD.n1098 AVDD.n1097 9.3005
R8452 AVDD.n1100 AVDD.n1099 9.3005
R8453 AVDD.n1103 AVDD.n1102 9.3005
R8454 AVDD.n1104 AVDD.n705 9.3005
R8455 AVDD.n1119 AVDD.n1118 9.3005
R8456 AVDD.n698 AVDD.n685 9.3005
R8457 AVDD.n1131 AVDD.n1129 9.3005
R8458 AVDD.n1141 AVDD.n573 9.3005
R8459 AVDD.n1141 AVDD.n572 9.3005
R8460 AVDD.n1141 AVDD.n574 9.3005
R8461 AVDD.n1141 AVDD.n571 9.3005
R8462 AVDD.n1141 AVDD.n575 9.3005
R8463 AVDD.n1141 AVDD.n570 9.3005
R8464 AVDD.n1141 AVDD.n576 9.3005
R8465 AVDD.n1141 AVDD.n569 9.3005
R8466 AVDD.n1141 AVDD.n577 9.3005
R8467 AVDD.n1141 AVDD.n568 9.3005
R8468 AVDD.n1141 AVDD.n578 9.3005
R8469 AVDD.n1141 AVDD.n567 9.3005
R8470 AVDD.n1141 AVDD.n579 9.3005
R8471 AVDD.n1141 AVDD.n566 9.3005
R8472 AVDD.n1141 AVDD.n580 9.3005
R8473 AVDD.n1141 AVDD.n565 9.3005
R8474 AVDD.n1141 AVDD.n581 9.3005
R8475 AVDD.n1141 AVDD.n564 9.3005
R8476 AVDD.n1118 AVDD.n1117 9.3005
R8477 AVDD.n698 AVDD.n697 9.3005
R8478 AVDD.n1132 AVDD.n1131 9.3005
R8479 AVDD.n1141 AVDD.n582 9.3005
R8480 AVDD.n1141 AVDD.n563 9.3005
R8481 AVDD.n1141 AVDD.n583 9.3005
R8482 AVDD.n1141 AVDD.n562 9.3005
R8483 AVDD.n1141 AVDD.n584 9.3005
R8484 AVDD.n1141 AVDD.n561 9.3005
R8485 AVDD.n1141 AVDD.n585 9.3005
R8486 AVDD.n1141 AVDD.n560 9.3005
R8487 AVDD.n1141 AVDD.n586 9.3005
R8488 AVDD.n1141 AVDD.n559 9.3005
R8489 AVDD.n1141 AVDD.n587 9.3005
R8490 AVDD.n1141 AVDD.n558 9.3005
R8491 AVDD.n1141 AVDD.n588 9.3005
R8492 AVDD.n1141 AVDD.n557 9.3005
R8493 AVDD.n1141 AVDD.n589 9.3005
R8494 AVDD.n1141 AVDD.n556 9.3005
R8495 AVDD.n1141 AVDD.n1140 9.3005
R8496 AVDD.n693 AVDD.n691 9.3005
R8497 AVDD.n1115 AVDD.n693 9.3005
R8498 AVDD.n1926 AVDD.n487 9.3005
R8499 AVDD.n1927 AVDD.n1926 9.3005
R8500 AVDD.n2849 AVDD.n2848 9.3005
R8501 AVDD.n450 AVDD.n448 9.3005
R8502 AVDD.n444 AVDD.n443 9.3005
R8503 AVDD.n2857 AVDD.n2856 9.3005
R8504 AVDD.n2859 AVDD.n2858 9.3005
R8505 AVDD.n438 AVDD.n435 9.3005
R8506 AVDD.n2866 AVDD.n2865 9.3005
R8507 AVDD.n436 AVDD.n432 9.3005
R8508 AVDD.n2871 AVDD.n2870 9.3005
R8509 AVDD.n406 AVDD.n405 9.3005
R8510 AVDD.n2903 AVDD.n2902 9.3005
R8511 AVDD.n2905 AVDD.n2904 9.3005
R8512 AVDD.n404 AVDD.n401 9.3005
R8513 AVDD.n403 AVDD.n397 9.3005
R8514 AVDD.n2913 AVDD.n2912 9.3005
R8515 AVDD.n2915 AVDD.n2914 9.3005
R8516 AVDD.n381 AVDD.n379 9.3005
R8517 AVDD.n375 AVDD.n374 9.3005
R8518 AVDD.n2945 AVDD.n2944 9.3005
R8519 AVDD.n351 AVDD.n343 9.3005
R8520 AVDD.n345 AVDD.n339 9.3005
R8521 AVDD.n2953 AVDD.n2952 9.3005
R8522 AVDD.n2955 AVDD.n2954 9.3005
R8523 AVDD.n337 AVDD.n335 9.3005
R8524 AVDD.n331 AVDD.n330 9.3005
R8525 AVDD.n2963 AVDD.n2962 9.3005
R8526 AVDD.n2965 AVDD.n2964 9.3005
R8527 AVDD.n308 AVDD.n302 9.3005
R8528 AVDD.n2995 AVDD.n2994 9.3005
R8529 AVDD.n2997 AVDD.n2996 9.3005
R8530 AVDD.n300 AVDD.n296 9.3005
R8531 AVDD.n299 AVDD.n291 9.3005
R8532 AVDD.n3005 AVDD.n3004 9.3005
R8533 AVDD.n3011 AVDD.n3010 9.3005
R8534 AVDD.n287 AVDD.n285 9.3005
R8535 AVDD.n281 AVDD.n280 9.3005
R8536 AVDD.n3042 AVDD.n3041 9.3005
R8537 AVDD.n258 AVDD.n255 9.3005
R8538 AVDD.n257 AVDD.n251 9.3005
R8539 AVDD.n3050 AVDD.n3049 9.3005
R8540 AVDD.n3056 AVDD.n3055 9.3005
R8541 AVDD.n247 AVDD.n245 9.3005
R8542 AVDD.n241 AVDD.n240 9.3005
R8543 AVDD.n3064 AVDD.n3063 9.3005
R8544 AVDD.n3066 AVDD.n3065 9.3005
R8545 AVDD.n217 AVDD.n212 9.3005
R8546 AVDD.n3096 AVDD.n3095 9.3005
R8547 AVDD.n3098 AVDD.n3097 9.3005
R8548 AVDD.n204 AVDD.n202 9.3005
R8549 AVDD.n197 AVDD.n196 9.3005
R8550 AVDD.n3106 AVDD.n3105 9.3005
R8551 AVDD.n3108 AVDD.n3107 9.3005
R8552 AVDD.n1730 AVDD.n195 9.3005
R8553 AVDD.n1728 AVDD.n1727 9.3005
R8554 AVDD.n1240 AVDD.n1230 9.3005
R8555 AVDD.n1233 AVDD.n1232 9.3005
R8556 AVDD.n1226 AVDD.n1225 9.3005
R8557 AVDD.n1751 AVDD.n1750 9.3005
R8558 AVDD.n1754 AVDD.n1753 9.3005
R8559 AVDD.n1198 AVDD.n1197 9.3005
R8560 AVDD.n1783 AVDD.n1782 9.3005
R8561 AVDD.n1785 AVDD.n1784 9.3005
R8562 AVDD.n1195 AVDD.n1193 9.3005
R8563 AVDD.n1189 AVDD.n1188 9.3005
R8564 AVDD.n1793 AVDD.n1792 9.3005
R8565 AVDD.n1795 AVDD.n1794 9.3005
R8566 AVDD.n1183 AVDD.n1180 9.3005
R8567 AVDD.n1802 AVDD.n1801 9.3005
R8568 AVDD.n1827 AVDD.n1826 9.3005
R8569 AVDD.n1155 AVDD.n1151 9.3005
R8570 AVDD.n1832 AVDD.n1831 9.3005
R8571 AVDD.n1149 AVDD.n1147 9.3005
R8572 AVDD.n1143 AVDD.n1142 9.3005
R8573 AVDD.n1840 AVDD.n1839 9.3005
R8574 AVDD.n1843 AVDD.n1842 9.3005
R8575 AVDD.n554 AVDD.n552 9.3005
R8576 AVDD.n548 AVDD.n547 9.3005
R8577 AVDD.n1874 AVDD.n1873 9.3005
R8578 AVDD.n526 AVDD.n523 9.3005
R8579 AVDD.n525 AVDD.n519 9.3005
R8580 AVDD.n1882 AVDD.n1881 9.3005
R8581 AVDD.n1888 AVDD.n1887 9.3005
R8582 AVDD.n515 AVDD.n512 9.3005
R8583 AVDD.n1895 AVDD.n1894 9.3005
R8584 AVDD.n1918 AVDD.n510 9.3005
R8585 AVDD.n1918 AVDD.n478 9.3005
R8586 AVDD.n1926 AVDD.n486 9.3005
R8587 AVDD.n1926 AVDD.n488 9.3005
R8588 AVDD.n1926 AVDD.n485 9.3005
R8589 AVDD.n1926 AVDD.n489 9.3005
R8590 AVDD.n1926 AVDD.n484 9.3005
R8591 AVDD.n1926 AVDD.n1925 9.3005
R8592 AVDD.n495 AVDD.n494 9.3005
R8593 AVDD.n493 AVDD.n492 9.3005
R8594 AVDD.n2840 AVDD.n2839 9.3005
R8595 AVDD.n453 AVDD.n451 9.3005
R8596 AVDD.n2847 AVDD.n2846 9.3005
R8597 AVDD.n430 AVDD.n427 9.3005
R8598 AVDD.n423 AVDD.n422 9.3005
R8599 AVDD.n2879 AVDD.n2878 9.3005
R8600 AVDD.n2881 AVDD.n2880 9.3005
R8601 AVDD.n421 AVDD.n418 9.3005
R8602 AVDD.n414 AVDD.n413 9.3005
R8603 AVDD.n2889 AVDD.n2888 9.3005
R8604 AVDD.n2895 AVDD.n2894 9.3005
R8605 AVDD.n2923 AVDD.n2922 9.3005
R8606 AVDD.n2925 AVDD.n2924 9.3005
R8607 AVDD.n367 AVDD.n365 9.3005
R8608 AVDD.n361 AVDD.n360 9.3005
R8609 AVDD.n2933 AVDD.n2932 9.3005
R8610 AVDD.n2936 AVDD.n2935 9.3005
R8611 AVDD.n355 AVDD.n353 9.3005
R8612 AVDD.n2943 AVDD.n2942 9.3005
R8613 AVDD.n328 AVDD.n326 9.3005
R8614 AVDD.n322 AVDD.n321 9.3005
R8615 AVDD.n2973 AVDD.n2972 9.3005
R8616 AVDD.n2975 AVDD.n2974 9.3005
R8617 AVDD.n316 AVDD.n313 9.3005
R8618 AVDD.n2982 AVDD.n2981 9.3005
R8619 AVDD.n314 AVDD.n310 9.3005
R8620 AVDD.n2987 AVDD.n2986 9.3005
R8621 AVDD.n3019 AVDD.n3018 9.3005
R8622 AVDD.n3021 AVDD.n3020 9.3005
R8623 AVDD.n274 AVDD.n271 9.3005
R8624 AVDD.n3028 AVDD.n3027 9.3005
R8625 AVDD.n272 AVDD.n268 9.3005
R8626 AVDD.n3033 AVDD.n3032 9.3005
R8627 AVDD.n266 AVDD.n261 9.3005
R8628 AVDD.n3040 AVDD.n3039 9.3005
R8629 AVDD.n234 AVDD.n231 9.3005
R8630 AVDD.n3073 AVDD.n3072 9.3005
R8631 AVDD.n232 AVDD.n228 9.3005
R8632 AVDD.n3078 AVDD.n3077 9.3005
R8633 AVDD.n226 AVDD.n223 9.3005
R8634 AVDD.n219 AVDD.n218 9.3005
R8635 AVDD.n3086 AVDD.n3085 9.3005
R8636 AVDD.n3088 AVDD.n3087 9.3005
R8637 AVDD.n1741 AVDD.n1740 9.3005
R8638 AVDD.n1743 AVDD.n1742 9.3005
R8639 AVDD.n1224 AVDD.n1222 9.3005
R8640 AVDD.n1218 AVDD.n1217 9.3005
R8641 AVDD.n1762 AVDD.n1761 9.3005
R8642 AVDD.n1765 AVDD.n1764 9.3005
R8643 AVDD.n1216 AVDD.n1208 9.3005
R8644 AVDD.n1210 AVDD.n1204 9.3005
R8645 AVDD.n1773 AVDD.n1772 9.3005
R8646 AVDD.n1775 AVDD.n1774 9.3005
R8647 AVDD.n1181 AVDD.n1177 9.3005
R8648 AVDD.n1807 AVDD.n1806 9.3005
R8649 AVDD.n1175 AVDD.n1172 9.3005
R8650 AVDD.n1168 AVDD.n1167 9.3005
R8651 AVDD.n1815 AVDD.n1814 9.3005
R8652 AVDD.n1817 AVDD.n1816 9.3005
R8653 AVDD.n1166 AVDD.n1163 9.3005
R8654 AVDD.n1160 AVDD.n1154 9.3005
R8655 AVDD.n1851 AVDD.n1850 9.3005
R8656 AVDD.n1853 AVDD.n1852 9.3005
R8657 AVDD.n542 AVDD.n539 9.3005
R8658 AVDD.n1860 AVDD.n1859 9.3005
R8659 AVDD.n540 AVDD.n536 9.3005
R8660 AVDD.n1865 AVDD.n1864 9.3005
R8661 AVDD.n534 AVDD.n529 9.3005
R8662 AVDD.n1872 AVDD.n1871 9.3005
R8663 AVDD.n1918 AVDD.n505 9.3005
R8664 AVDD.n1919 AVDD.n1918 9.3005
R8665 AVDD.n1918 AVDD.n508 9.3005
R8666 AVDD.n1918 AVDD.n1896 9.3005
R8667 AVDD.n1918 AVDD.n507 9.3005
R8668 AVDD.n1918 AVDD.n1917 9.3005
R8669 AVDD.n1928 AVDD.n464 9.3005
R8670 AVDD.n2834 AVDD.n2833 9.3005
R8671 AVDD.n2388 AVDD.n468 9.3005
R8672 AVDD.n2393 AVDD.n2392 9.3005
R8673 AVDD.n2390 AVDD.n2385 9.3005
R8674 AVDD.n2398 AVDD.n2397 9.3005
R8675 AVDD.n2411 AVDD.n2410 9.3005
R8676 AVDD.n2439 AVDD.n2438 9.3005
R8677 AVDD.n2443 AVDD.n2442 9.3005
R8678 AVDD.n2449 AVDD.n2448 9.3005
R8679 AVDD.n2451 AVDD.n2369 9.3005
R8680 AVDD.n2520 AVDD.n2519 9.3005
R8681 AVDD.n2516 AVDD.n2515 9.3005
R8682 AVDD.n2456 AVDD.n2454 9.3005
R8683 AVDD.n2511 AVDD.n2510 9.3005
R8684 AVDD.n2508 AVDD.n2507 9.3005
R8685 AVDD.n2485 AVDD.n2484 9.3005
R8686 AVDD.n2527 AVDD.n2526 9.3005
R8687 AVDD.n2535 AVDD.n2534 9.3005
R8688 AVDD.n2532 AVDD.n2531 9.3005
R8689 AVDD.n2541 AVDD.n2540 9.3005
R8690 AVDD.n2544 AVDD.n2359 9.3005
R8691 AVDD.n2549 AVDD.n2548 9.3005
R8692 AVDD.n2546 AVDD.n2358 9.3005
R8693 AVDD.n2554 AVDD.n2553 9.3005
R8694 AVDD.n2592 AVDD.n2591 9.3005
R8695 AVDD.n2595 AVDD.n2343 9.3005
R8696 AVDD.n2601 AVDD.n2600 9.3005
R8697 AVDD.n2598 AVDD.n2597 9.3005
R8698 AVDD.n2607 AVDD.n2606 9.3005
R8699 AVDD.n2610 AVDD.n2340 9.3005
R8700 AVDD.n2615 AVDD.n2614 9.3005
R8701 AVDD.n2612 AVDD.n2339 9.3005
R8702 AVDD.n2620 AVDD.n2619 9.3005
R8703 AVDD.n2633 AVDD.n2632 9.3005
R8704 AVDD.n2626 AVDD.n2625 9.3005
R8705 AVDD.n2587 AVDD.n2586 9.3005
R8706 AVDD.n2584 AVDD.n2347 9.3005
R8707 AVDD.n2582 AVDD.n2581 9.3005
R8708 AVDD.n2571 AVDD.n2570 9.3005
R8709 AVDD.n2566 AVDD.n2351 9.3005
R8710 AVDD.n2564 AVDD.n2350 9.3005
R8711 AVDD.n2562 AVDD.n2561 9.3005
R8712 AVDD.n2560 AVDD.n2559 9.3005
R8713 AVDD.n2488 AVDD.n2487 9.3005
R8714 AVDD.n2490 AVDD.n2489 9.3005
R8715 AVDD.n2493 AVDD.n2492 9.3005
R8716 AVDD.n2478 AVDD.n2473 9.3005
R8717 AVDD.n2498 AVDD.n2497 9.3005
R8718 AVDD.n2500 AVDD.n2460 9.3005
R8719 AVDD.n2503 AVDD.n2502 9.3005
R8720 AVDD.n2461 AVDD.n2459 9.3005
R8721 AVDD.n2435 AVDD.n2434 9.3005
R8722 AVDD.n2432 AVDD.n2374 9.3005
R8723 AVDD.n2430 AVDD.n2429 9.3005
R8724 AVDD.n2421 AVDD.n2420 9.3005
R8725 AVDD.n2424 AVDD.n2423 9.3005
R8726 AVDD.n2418 AVDD.n2378 9.3005
R8727 AVDD.n2416 AVDD.n2415 9.3005
R8728 AVDD.n2400 AVDD.n2382 9.3005
R8729 AVDD.n3108 AVDD.n194 8.65932
R8730 AVDD.n3110 AVDD.n3109 8.65932
R8731 AVDD.n975 AVDD.n974 8.65932
R8732 AVDD.n1102 AVDD.n1101 8.65932
R8733 AVDD.n981 AVDD.n979 8.65932
R8734 AVDD.n723 AVDD.n710 8.65932
R8735 AVDD.n3105 AVDD.n3104 8.28285
R8736 AVDD.n232 AVDD.n224 8.28285
R8737 AVDD.n3057 AVDD.n245 8.28285
R8738 AVDD.n3026 AVDD.n274 8.28285
R8739 AVDD.n3004 AVDD.n3003 8.28285
R8740 AVDD.n2972 AVDD.n320 8.28285
R8741 AVDD.n2956 AVDD.n335 8.28285
R8742 AVDD.n365 AVDD.n363 8.28285
R8743 AVDD.n2912 AVDD.n2911 8.28285
R8744 AVDD.n2878 AVDD.n419 8.28285
R8745 AVDD.n2860 AVDD.n438 8.28285
R8746 AVDD.n1335 AVDD.n1334 8.28285
R8747 AVDD.n1379 AVDD.n1376 8.28285
R8748 AVDD.n1692 AVDD.n1691 8.28285
R8749 AVDD.n1649 AVDD.n1402 8.28285
R8750 AVDD.n1626 AVDD.n1625 8.28285
R8751 AVDD.n1596 AVDD.n1461 8.28285
R8752 AVDD.n1574 AVDD.n1491 8.28285
R8753 AVDD.n1538 AVDD.n1506 8.28285
R8754 AVDD.n1517 AVDD.n9 8.28285
R8755 AVDD.n2271 AVDD.n2270 8.28285
R8756 AVDD.n2297 AVDD.n2222 8.28285
R8757 AVDD.n1902 AVDD.n485 8.28285
R8758 AVDD.n2833 AVDD.n2832 8.28285
R8759 AVDD.n2430 AVDD.n2376 8.28285
R8760 AVDD.n2452 AVDD.n2451 8.28285
R8761 AVDD.n2492 AVDD.n2480 8.28285
R8762 AVDD.n2532 AVDD.n2360 8.28285
R8763 AVDD.n2582 AVDD.n2348 8.28285
R8764 AVDD.n2598 AVDD.n2341 8.28285
R8765 AVDD.n2209 AVDD.n2190 8.28285
R8766 AVDD.n1889 AVDD.n512 8.28285
R8767 AVDD.n1858 AVDD.n542 8.28285
R8768 AVDD.n1839 AVDD.n1838 8.28285
R8769 AVDD.n1172 AVDD.n1170 8.28285
R8770 AVDD.n1792 AVDD.n1791 8.28285
R8771 AVDD.n1761 AVDD.n1209 8.28285
R8772 AVDD.n1905 AVDD.n1896 8.28285
R8773 AVDD.n2828 AVDD.n475 8.28285
R8774 AVDD.n2797 AVDD.n1968 8.28285
R8775 AVDD.n2778 AVDD.n1999 8.28285
R8776 AVDD.n2746 AVDD.n2032 8.28285
R8777 AVDD.n2726 AVDD.n2058 8.28285
R8778 AVDD.n2695 AVDD.n2106 8.28285
R8779 AVDD.n2675 AVDD.n2131 8.28285
R8780 AVDD.n2205 AVDD.n2177 8.28285
R8781 AVDD.n3293 AVDD.n99 8.28285
R8782 AVDD.n3256 AVDD.n113 8.28285
R8783 AVDD.n3237 AVDD.n3236 8.28285
R8784 AVDD.n3204 AVDD.n145 8.28285
R8785 AVDD.n3186 AVDD.n3185 8.28285
R8786 AVDD.n3146 AVDD.n171 8.28285
R8787 AVDD.n948 AVDD.n784 8.28285
R8788 AVDD.n911 AVDD.n806 8.28285
R8789 AVDD.n892 AVDD.n891 8.28285
R8790 AVDD.n856 AVDD.n855 8.28285
R8791 AVDD.n601 AVDD.n580 8.28285
R8792 AVDD.n628 AVDD.n560 8.28285
R8793 AVDD.n646 AVDD.n570 8.28285
R8794 AVDD.n673 AVDD.n556 8.28285
R8795 AVDD.n1024 AVDD.n752 7.90638
R8796 AVDD.n1017 AVDD.n759 7.90638
R8797 AVDD.n1100 AVDD.n716 7.15344
R8798 AVDD.n1091 AVDD.n1090 7.15344
R8799 AVDD.n777 AVDD.t130 6.92038
R8800 AVDD.n199 AVDD.n197 6.77697
R8801 AVDD.n3079 AVDD.n3078 6.77697
R8802 AVDD.n3056 AVDD.n246 6.77697
R8803 AVDD.n3027 AVDD.n273 6.77697
R8804 AVDD.n293 AVDD.n291 6.77697
R8805 AVDD.n2976 AVDD.n2975 6.77697
R8806 AVDD.n2955 AVDD.n336 6.77697
R8807 AVDD.n2931 AVDD.n361 6.77697
R8808 AVDD.n399 AVDD.n397 6.77697
R8809 AVDD.n2882 AVDD.n2881 6.77697
R8810 AVDD.n2859 AVDD.n442 6.77697
R8811 AVDD.n496 AVDD.n495 6.77697
R8812 AVDD.n1346 AVDD.n1345 6.77697
R8813 AVDD.n1380 AVDD.n1375 6.77697
R8814 AVDD.n1688 AVDD.n1394 6.77697
R8815 AVDD.n1653 AVDD.n1652 6.77697
R8816 AVDD.n1622 AVDD.n1444 6.77697
R8817 AVDD.n1600 AVDD.n1597 6.77697
R8818 AVDD.n1573 AVDD.n1492 6.77697
R8819 AVDD.n1542 AVDD.n1539 6.77697
R8820 AVDD.n3301 AVDD.n3300 6.77697
R8821 AVDD.n2267 AVDD.n2266 6.77697
R8822 AVDD.n2302 AVDD.n2301 6.77697
R8823 AVDD.n2322 AVDD.n2321 6.77697
R8824 AVDD.n499 AVDD.n489 6.77697
R8825 AVDD.n2389 AVDD.n468 6.77697
R8826 AVDD.n2422 AVDD.n2421 6.77697
R8827 AVDD.n2519 AVDD.n2518 6.77697
R8828 AVDD.n2478 AVDD.n2471 6.77697
R8829 AVDD.n2543 AVDD.n2541 6.77697
R8830 AVDD.n2570 AVDD.n2569 6.77697
R8831 AVDD.n2609 AVDD.n2607 6.77697
R8832 AVDD.n2210 AVDD.n2196 6.77697
R8833 AVDD.n1888 AVDD.n514 6.77697
R8834 AVDD.n1859 AVDD.n541 6.77697
R8835 AVDD.n1145 AVDD.n1143 6.77697
R8836 AVDD.n1813 AVDD.n1168 6.77697
R8837 AVDD.n1191 AVDD.n1189 6.77697
R8838 AVDD.n1766 AVDD.n1765 6.77697
R8839 AVDD.n508 AVDD.n506 6.77697
R8840 AVDD.n2827 AVDD.n476 6.77697
R8841 AVDD.n2803 AVDD.n2802 6.77697
R8842 AVDD.n2777 AVDD.n2000 6.77697
R8843 AVDD.n2752 AVDD.n2751 6.77697
R8844 AVDD.n2725 AVDD.n2059 6.77697
R8845 AVDD.n2105 AVDD.n2100 6.77697
R8846 AVDD.n2674 AVDD.n2132 6.77697
R8847 AVDD.n2171 AVDD.n2169 6.77697
R8848 AVDD.n107 AVDD.n106 6.77697
R8849 AVDD.n3260 AVDD.n3259 6.77697
R8850 AVDD.n3233 AVDD.n3232 6.77697
R8851 AVDD.n3208 AVDD.n3205 6.77697
R8852 AVDD.n3182 AVDD.n3181 6.77697
R8853 AVDD.n3150 AVDD.n3147 6.77697
R8854 AVDD.n947 AVDD.n786 6.77697
R8855 AVDD.n915 AVDD.n914 6.77697
R8856 AVDD.n887 AVDD.n822 6.77697
R8857 AVDD.n860 AVDD.n843 6.77697
R8858 AVDD.n603 AVDD.n566 6.77697
R8859 AVDD.n626 AVDD.n585 6.77697
R8860 AVDD.n648 AVDD.n575 6.77697
R8861 AVDD.n671 AVDD.n589 6.77697
R8862 AVDD.n1032 AVDD.n1030 6.4005
R8863 AVDD.n1007 AVDD.n750 6.4005
R8864 AVDD.n1097 AVDD.n1096 5.64756
R8865 AVDD.n727 AVDD.n722 5.64756
R8866 AVDD.t0 AVDD.n1060 5.6023
R8867 AVDD.n1922 AVDD.n501 5.56371
R8868 AVDD.n1922 AVDD.n502 5.56371
R8869 AVDD.n1909 AVDD.n1904 5.56371
R8870 AVDD.n1910 AVDD.n1909 5.56371
R8871 AVDD.n1914 AVDD.n480 5.56371
R8872 AVDD.n1931 AVDD.n480 5.56371
R8873 AVDD.n1931 AVDD.n471 5.56371
R8874 AVDD.n2830 AVDD.n471 5.56371
R8875 AVDD.n2830 AVDD.n472 5.56371
R8876 AVDD.n2821 AVDD.n472 5.56371
R8877 AVDD.n2820 AVDD.n2819 5.56371
R8878 AVDD.n2819 AVDD.n1945 5.56371
R8879 AVDD.n2406 AVDD.n1945 5.56371
R8880 AVDD.n2807 AVDD.n1961 5.56371
R8881 AVDD.n2807 AVDD.n2806 5.56371
R8882 AVDD.n2806 AVDD.n2805 5.56371
R8883 AVDD.n2794 AVDD.n1978 5.56371
R8884 AVDD.n2794 AVDD.n2793 5.56371
R8885 AVDD.n2793 AVDD.t16 5.56371
R8886 AVDD.t16 AVDD.n1981 5.56371
R8887 AVDD.n2782 AVDD.n1981 5.56371
R8888 AVDD.n2782 AVDD.n2781 5.56371
R8889 AVDD.n2781 AVDD.n2780 5.56371
R8890 AVDD.n2780 AVDD.n1996 5.56371
R8891 AVDD.n2770 AVDD.n1996 5.56371
R8892 AVDD.n2769 AVDD.n2768 5.56371
R8893 AVDD.n2768 AVDD.n2009 5.56371
R8894 AVDD.n2467 AVDD.n2009 5.56371
R8895 AVDD.n2756 AVDD.n2025 5.56371
R8896 AVDD.n2756 AVDD.n2755 5.56371
R8897 AVDD.n2755 AVDD.n2754 5.56371
R8898 AVDD.n2743 AVDD.n2037 5.56371
R8899 AVDD.n2743 AVDD.n2742 5.56371
R8900 AVDD.n2742 AVDD.n2741 5.56371
R8901 AVDD.n2730 AVDD.n2051 5.56371
R8902 AVDD.n2730 AVDD.n2729 5.56371
R8903 AVDD.n2728 AVDD.n2055 5.56371
R8904 AVDD.n2718 AVDD.n2055 5.56371
R8905 AVDD.n2718 AVDD.n2717 5.56371
R8906 AVDD.n2716 AVDD.n2078 5.56371
R8907 AVDD.n2092 AVDD.n2078 5.56371
R8908 AVDD.n2706 AVDD.n2092 5.56371
R8909 AVDD.n2706 AVDD.n2705 5.56371
R8910 AVDD.n2705 AVDD.n2704 5.56371
R8911 AVDD.n2704 AVDD.n2096 5.56371
R8912 AVDD.n2692 AVDD.n2110 5.56371
R8913 AVDD.n2692 AVDD.n2691 5.56371
R8914 AVDD.n2691 AVDD.n2690 5.56371
R8915 AVDD.n2679 AVDD.n2124 5.56371
R8916 AVDD.n2679 AVDD.n2678 5.56371
R8917 AVDD.n2677 AVDD.n2128 5.56371
R8918 AVDD.n2667 AVDD.n2128 5.56371
R8919 AVDD.n2667 AVDD.n2666 5.56371
R8920 AVDD.n2665 AVDD.n2147 5.56371
R8921 AVDD.n2161 AVDD.n2147 5.56371
R8922 AVDD.n2655 AVDD.n2161 5.56371
R8923 AVDD.n2655 AVDD.n2654 5.56371
R8924 AVDD.n2654 AVDD.n2653 5.56371
R8925 AVDD.n2653 AVDD.n2165 5.56371
R8926 AVDD.n2207 AVDD.n2202 5.56371
R8927 AVDD.n2202 AVDD.n2182 5.56371
R8928 AVDD.n2645 AVDD.n2182 5.56371
R8929 AVDD.n2644 AVDD.n2643 5.56371
R8930 AVDD.n2643 AVDD.n13 5.56371
R8931 AVDD.n1910 AVDD.t134 5.4819
R8932 AVDD.n2051 AVDD.t32 5.40009
R8933 AVDD.n3099 AVDD.n202 5.27109
R8934 AVDD.n223 AVDD.n221 5.27109
R8935 AVDD.n3049 AVDD.n3048 5.27109
R8936 AVDD.n272 AVDD.n265 5.27109
R8937 AVDD.n2998 AVDD.n296 5.27109
R8938 AVDD.n2980 AVDD.n316 5.27109
R8939 AVDD.n2952 AVDD.n2951 5.27109
R8940 AVDD.n2932 AVDD.n359 5.27109
R8941 AVDD.n2906 AVDD.n401 5.27109
R8942 AVDD.n418 AVDD.n416 5.27109
R8943 AVDD.n2856 AVDD.n2855 5.27109
R8944 AVDD.n492 AVDD.n457 5.27109
R8945 AVDD.n1349 AVDD.n1332 5.27109
R8946 AVDD.n1372 AVDD.n1327 5.27109
R8947 AVDD.n1681 AVDD.n1680 5.27109
R8948 AVDD.n1656 AVDD.n1401 5.27109
R8949 AVDD.n1619 AVDD.n1618 5.27109
R8950 AVDD.n1601 AVDD.n1453 5.27109
R8951 AVDD.n1570 AVDD.n1569 5.27109
R8952 AVDD.n1543 AVDD.n1504 5.27109
R8953 AVDD.n2235 AVDD.n10 5.27109
R8954 AVDD.n2263 AVDD.n2229 5.27109
R8955 AVDD.n2305 AVDD.n2221 5.27109
R8956 AVDD.n2325 AVDD.n2323 5.27109
R8957 AVDD.n1924 AVDD.n484 5.27109
R8958 AVDD.n2392 AVDD.n2391 5.27109
R8959 AVDD.n2423 AVDD.n2419 5.27109
R8960 AVDD.n2516 AVDD.n2453 5.27109
R8961 AVDD.n2499 AVDD.n2498 5.27109
R8962 AVDD.n2545 AVDD.n2544 5.27109
R8963 AVDD.n2566 AVDD.n2565 5.27109
R8964 AVDD.n2611 AVDD.n2610 5.27109
R8965 AVDD.n2635 AVDD.n2189 5.27109
R8966 AVDD.n1881 AVDD.n1880 5.27109
R8967 AVDD.n540 AVDD.n533 5.27109
R8968 AVDD.n1833 AVDD.n1147 5.27109
R8969 AVDD.n1814 AVDD.n1164 5.27109
R8970 AVDD.n1786 AVDD.n1193 5.27109
R8971 AVDD.n1208 AVDD.n1206 5.27109
R8972 AVDD.n1920 AVDD.n1919 5.27109
R8973 AVDD.n2824 AVDD.n2823 5.27109
R8974 AVDD.n1967 AVDD.n1966 5.27109
R8975 AVDD.n2773 AVDD.n2772 5.27109
R8976 AVDD.n2031 AVDD.n2030 5.27109
R8977 AVDD.n2721 AVDD.n2720 5.27109
R8978 AVDD.n2702 AVDD.n2701 5.27109
R8979 AVDD.n2670 AVDD.n2669 5.27109
R8980 AVDD.n2651 AVDD.n2650 5.27109
R8981 AVDD.n3287 AVDD.n3286 5.27109
R8982 AVDD.n3263 AVDD.n112 5.27109
R8983 AVDD.n3229 AVDD.n128 5.27109
R8984 AVDD.n3209 AVDD.n141 5.27109
R8985 AVDD.n3178 AVDD.n161 5.27109
R8986 AVDD.n3151 AVDD.n168 5.27109
R8987 AVDD.n942 AVDD.n941 5.27109
R8988 AVDD.n919 AVDD.n804 5.27109
R8989 AVDD.n886 AVDD.n825 5.27109
R8990 AVDD.n861 AVDD.n840 5.27109
R8991 AVDD.n606 AVDD.n579 5.27109
R8992 AVDD.n623 AVDD.n561 5.27109
R8993 AVDD.n651 AVDD.n571 5.27109
R8994 AVDD.n668 AVDD.n557 5.27109
R8995 AVDD.n2124 AVDD.t29 5.23646
R8996 AVDD.t192 AVDD.n2644 5.07284
R8997 AVDD.n1031 AVDD.n737 4.89462
R8998 AVDD.n1037 AVDD.n748 4.89462
R8999 AVDD.n2678 AVDD.t18 4.74559
R9000 AVDD.n2837 AVDD.n2836 4.61479
R9001 AVDD.n2729 AVDD.t35 4.58197
R9002 AVDD.n1267 AVDD.n1248 4.53153
R9003 AVDD.n1292 AVDD.n1273 4.53153
R9004 AVDD.n1713 AVDD.n190 4.53153
R9005 AVDD.n1703 AVDD.n1299 4.53153
R9006 AVDD.n1433 AVDD.n1432 4.53153
R9007 AVDD.n1487 AVDD.n1486 4.53153
R9008 AVDD.n3304 AVDD.n2 4.53153
R9009 AVDD.n2631 AVDD.n2630 4.53153
R9010 AVDD.n1259 AVDD.n1258 4.5005
R9011 AVDD.n1256 AVDD.n1250 4.5005
R9012 AVDD.n1255 AVDD.n1254 4.5005
R9013 AVDD.n1270 AVDD.n1269 4.5005
R9014 AVDD.n1268 AVDD.n1265 4.5005
R9015 AVDD.n1284 AVDD.n1283 4.5005
R9016 AVDD.n1281 AVDD.n1275 4.5005
R9017 AVDD.n1280 AVDD.n1279 4.5005
R9018 AVDD.n1295 AVDD.n1294 4.5005
R9019 AVDD.n1293 AVDD.n1290 4.5005
R9020 AVDD.n1720 AVDD.n1719 4.5005
R9021 AVDD.n1721 AVDD.n1241 4.5005
R9022 AVDD.n1723 AVDD.n1722 4.5005
R9023 AVDD.n1710 AVDD.n1247 4.5005
R9024 AVDD.n1712 AVDD.n1711 4.5005
R9025 AVDD.n1310 AVDD.n1309 4.5005
R9026 AVDD.n1307 AVDD.n1301 4.5005
R9027 AVDD.n1306 AVDD.n1305 4.5005
R9028 AVDD.n1706 AVDD.n1705 4.5005
R9029 AVDD.n1704 AVDD.n1316 4.5005
R9030 AVDD.n1421 AVDD.n1420 4.5005
R9031 AVDD.n1418 AVDD.n1412 4.5005
R9032 AVDD.n1417 AVDD.n1416 4.5005
R9033 AVDD.n1430 AVDD.n1429 4.5005
R9034 AVDD.n1431 AVDD.n1410 4.5005
R9035 AVDD.n1475 AVDD.n1474 4.5005
R9036 AVDD.n1472 AVDD.n1466 4.5005
R9037 AVDD.n1471 AVDD.n1470 4.5005
R9038 AVDD.n1484 AVDD.n1483 4.5005
R9039 AVDD.n1485 AVDD.n1464 4.5005
R9040 AVDD.n391 AVDD.n390 4.5005
R9041 AVDD.n392 AVDD.n383 4.5005
R9042 AVDD.n394 AVDD.n393 4.5005
R9043 AVDD.n3307 AVDD.n3306 4.5005
R9044 AVDD.n3305 AVDD.n5 4.5005
R9045 AVDD.n2354 AVDD.n2353 4.5005
R9046 AVDD.n2575 AVDD.n2574 4.5005
R9047 AVDD.n2577 AVDD.n2576 4.5005
R9048 AVDD.n2364 AVDD.n2352 4.5005
R9049 AVDD.n2523 AVDD.n2363 4.5005
R9050 AVDD.n2525 AVDD.n2524 4.5005
R9051 AVDD.n2522 AVDD.n2521 4.5005
R9052 AVDD.n2447 AVDD.n2368 4.5005
R9053 AVDD.n2446 AVDD.n2445 4.5005
R9054 AVDD.n466 AVDD.n465 4.5005
R9055 AVDD.n2836 AVDD.n2835 4.5005
R9056 AVDD.n2629 AVDD.n2212 4.5005
R9057 AVDD.n2628 AVDD.n2627 4.5005
R9058 AVDD.n1904 AVDD.t141 4.50016
R9059 AVDD.n1978 AVDD.t23 4.41834
R9060 AVDD.n1123 AVDD.t149 4.28423
R9061 AVDD.n2037 AVDD.t15 4.25472
R9062 AVDD.n3108 AVDD.n193 4.14168
R9063 AVDD.n3109 AVDD.n192 4.14168
R9064 AVDD.n733 AVDD.n718 4.14168
R9065 AVDD.n1081 AVDD.n728 4.14168
R9066 AVDD.n2110 AVDD.t8 4.0911
R9067 AVDD.n2207 AVDD.t144 3.92747
R9068 AVDD.n3098 AVDD.n203 3.76521
R9069 AVDD.n3084 AVDD.n219 3.76521
R9070 AVDD.n253 AVDD.n251 3.76521
R9071 AVDD.n3034 AVDD.n3033 3.76521
R9072 AVDD.n2981 AVDD.n315 3.76521
R9073 AVDD.n341 AVDD.n339 3.76521
R9074 AVDD.n2937 AVDD.n2936 3.76521
R9075 AVDD.n2905 AVDD.n402 3.76521
R9076 AVDD.n2887 AVDD.n414 3.76521
R9077 AVDD.n446 AVDD.n444 3.76521
R9078 AVDD.n2841 AVDD.n2840 3.76521
R9079 AVDD.n1353 AVDD.n1350 3.76521
R9080 AVDD.n1371 AVDD.n1328 3.76521
R9081 AVDD.n1677 AVDD.n1397 3.76521
R9082 AVDD.n1660 AVDD.n1657 3.76521
R9083 AVDD.n1605 AVDD.n1604 3.76521
R9084 AVDD.n1566 AVDD.n1495 3.76521
R9085 AVDD.n1548 AVDD.n1547 3.76521
R9086 AVDD.n2238 AVDD.n2237 3.76521
R9087 AVDD.n2262 AVDD.n2230 3.76521
R9088 AVDD.n2309 AVDD.n2306 3.76521
R9089 AVDD.n2329 AVDD.n2326 3.76521
R9090 AVDD.n1925 AVDD.n490 3.76521
R9091 AVDD.n2390 AVDD.n2384 3.76521
R9092 AVDD.n2418 AVDD.n2417 3.76521
R9093 AVDD.n2457 AVDD.n2456 3.76521
R9094 AVDD.n2501 AVDD.n2500 3.76521
R9095 AVDD.n2548 AVDD.n2547 3.76521
R9096 AVDD.n2564 AVDD.n2563 3.76521
R9097 AVDD.n2614 AVDD.n2613 3.76521
R9098 AVDD.n2636 AVDD.n2634 3.76521
R9099 AVDD.n521 AVDD.n519 3.76521
R9100 AVDD.n1866 AVDD.n1865 3.76521
R9101 AVDD.n1832 AVDD.n1148 3.76521
R9102 AVDD.n1818 AVDD.n1817 3.76521
R9103 AVDD.n1785 AVDD.n1194 3.76521
R9104 AVDD.n1771 AVDD.n1204 3.76521
R9105 AVDD.n511 AVDD.n505 3.76521
R9106 AVDD.n1947 AVDD.n1940 3.76521
R9107 AVDD.n2809 AVDD.n1958 3.76521
R9108 AVDD.n2011 AVDD.n2004 3.76521
R9109 AVDD.n2758 AVDD.n2022 3.76521
R9110 AVDD.n2080 AVDD.n2073 3.76521
R9111 AVDD.n2099 AVDD.n2098 3.76521
R9112 AVDD.n2149 AVDD.n2142 3.76521
R9113 AVDD.n2168 AVDD.n2167 3.76521
R9114 AVDD.n3284 AVDD.n108 3.76521
R9115 AVDD.n3267 AVDD.n3264 3.76521
R9116 AVDD.n3228 AVDD.n129 3.76521
R9117 AVDD.n3213 AVDD.n3212 3.76521
R9118 AVDD.n3177 AVDD.n162 3.76521
R9119 AVDD.n3161 AVDD.n3158 3.76521
R9120 AVDD.n937 AVDD.n790 3.76521
R9121 AVDD.n920 AVDD.n799 3.76521
R9122 AVDD.n883 AVDD.n882 3.76521
R9123 AVDD.n865 AVDD.n864 3.76521
R9124 AVDD.n608 AVDD.n567 3.76521
R9125 AVDD.n621 AVDD.n584 3.76521
R9126 AVDD.n653 AVDD.n574 3.76521
R9127 AVDD.n666 AVDD.n588 3.76521
R9128 AVDD.n2770 AVDD.t11 3.60022
R9129 AVDD.n2666 AVDD.t38 3.60022
R9130 AVDD.n1254 AVDD.n1253 3.47788
R9131 AVDD.n1279 AVDD.n1278 3.47788
R9132 AVDD.n1725 AVDD.n1723 3.47788
R9133 AVDD.n1305 AVDD.n1304 3.47788
R9134 AVDD.n1470 AVDD.n1469 3.47788
R9135 AVDD.n395 AVDD.n394 3.47788
R9136 AVDD.n1416 AVDD.n1415 3.47615
R9137 AVDD.n2821 AVDD.t20 3.4366
R9138 AVDD.n2717 AVDD.t19 3.4366
R9139 AVDD.n2336 AVDD.n1 3.4105
R9140 AVDD.n3309 AVDD.n3308 3.4105
R9141 AVDD.n1481 AVDD.n0 3.4105
R9142 AVDD.n1427 AVDD.n1298 3.4105
R9143 AVDD.n1708 AVDD.n1707 3.4105
R9144 AVDD.n1715 AVDD.n1714 3.4105
R9145 AVDD.n1297 AVDD.n1296 3.4105
R9146 AVDD.n1272 AVDD.n1271 3.4105
R9147 AVDD.n1065 AVDD.n1064 3.38874
R9148 AVDD.n1039 AVDD.n1038 3.38874
R9149 AVDD.t27 AVDD.n1961 3.27298
R9150 AVDD.t22 AVDD.n2025 3.10935
R9151 AVDD.n2997 AVDD.n297 2.63579
R9152 AVDD.n1446 AVDD.n298 2.63579
R9153 AVDD.n1076 AVDD.n1075 2.63579
R9154 AVDD.n1082 AVDD.n726 2.63579
R9155 AVDD.n2467 AVDD.t22 2.45486
R9156 AVDD.n2406 AVDD.t27 2.29123
R9157 AVDD.n3095 AVDD.n3094 2.25932
R9158 AVDD.n3085 AVDD.n216 2.25932
R9159 AVDD.n3043 AVDD.n255 2.25932
R9160 AVDD.n3038 AVDD.n261 2.25932
R9161 AVDD.n2994 AVDD.n2993 2.25932
R9162 AVDD.n314 AVDD.n307 2.25932
R9163 AVDD.n2946 AVDD.n343 2.25932
R9164 AVDD.n2941 AVDD.n355 2.25932
R9165 AVDD.n2902 AVDD.n2901 2.25932
R9166 AVDD.n2888 AVDD.n410 2.25932
R9167 AVDD.n2850 AVDD.n448 2.25932
R9168 AVDD.n2845 AVDD.n453 2.25932
R9169 AVDD.n1354 AVDD.n1330 2.25932
R9170 AVDD.n1367 AVDD.n1366 2.25932
R9171 AVDD.n1674 AVDD.n1673 2.25932
R9172 AVDD.n1661 AVDD.n1399 2.25932
R9173 AVDD.n1615 AVDD.n1614 2.25932
R9174 AVDD.n1608 AVDD.n1452 2.25932
R9175 AVDD.n1559 AVDD.n1558 2.25932
R9176 AVDD.n1551 AVDD.n1503 2.25932
R9177 AVDD.n2241 AVDD.n2234 2.25932
R9178 AVDD.n2257 AVDD.n2256 2.25932
R9179 AVDD.n2310 AVDD.n2219 2.25932
R9180 AVDD.n2330 AVDD.n2319 2.25932
R9181 AVDD.n2399 AVDD.n2398 2.25932
R9182 AVDD.n2416 AVDD.n2381 2.25932
R9183 AVDD.n2510 AVDD.n2509 2.25932
R9184 AVDD.n2502 AVDD.n2470 2.25932
R9185 AVDD.n2546 AVDD.n2357 2.25932
R9186 AVDD.n2562 AVDD.n2355 2.25932
R9187 AVDD.n2612 AVDD.n2338 2.25932
R9188 AVDD.n2633 AVDD.n2211 2.25932
R9189 AVDD.n1875 AVDD.n523 2.25932
R9190 AVDD.n1870 AVDD.n529 2.25932
R9191 AVDD.n1156 AVDD.n1155 2.25932
R9192 AVDD.n1163 AVDD.n1161 2.25932
R9193 AVDD.n1782 AVDD.n1781 2.25932
R9194 AVDD.n1772 AVDD.n1202 2.25932
R9195 AVDD.n2817 AVDD.n1948 2.25932
R9196 AVDD.n2810 AVDD.n1957 2.25932
R9197 AVDD.n2766 AVDD.n2012 2.25932
R9198 AVDD.n2759 AVDD.n2021 2.25932
R9199 AVDD.n2714 AVDD.n2081 2.25932
R9200 AVDD.n2708 AVDD.n2089 2.25932
R9201 AVDD.n2663 AVDD.n2150 2.25932
R9202 AVDD.n2657 AVDD.n2158 2.25932
R9203 AVDD.n3281 AVDD.n3280 2.25932
R9204 AVDD.n3268 AVDD.n110 2.25932
R9205 AVDD.n139 AVDD.n136 2.25932
R9206 AVDD.n3216 AVDD.n140 2.25932
R9207 AVDD.n3174 AVDD.n3173 2.25932
R9208 AVDD.n3162 AVDD.n166 2.25932
R9209 AVDD.n936 AVDD.n793 2.25932
R9210 AVDD.n926 AVDD.n925 2.25932
R9211 AVDD.n878 AVDD.n831 2.25932
R9212 AVDD.n871 AVDD.n838 2.25932
R9213 AVDD.n612 AVDD.n578 2.25932
R9214 AVDD.n618 AVDD.n562 2.25932
R9215 AVDD.n657 AVDD.n572 2.25932
R9216 AVDD.n663 AVDD.n558 2.25932
R9217 AVDD.t20 AVDD.n2820 2.12761
R9218 AVDD.t19 AVDD.n2716 2.12761
R9219 AVDD.n2445 AVDD.n465 1.96479
R9220 AVDD.t11 AVDD.n2769 1.96399
R9221 AVDD.t38 AVDD.n2665 1.96399
R9222 AVDD.n1051 AVDD.n738 1.88285
R9223 AVDD.n1041 AVDD.n1040 1.88285
R9224 AVDD.n1263 AVDD.n1259 1.87264
R9225 AVDD.n1288 AVDD.n1284 1.87264
R9226 AVDD.n1719 AVDD.n1718 1.87264
R9227 AVDD.n1314 AVDD.n1310 1.87264
R9228 AVDD.n1479 AVDD.n1475 1.87264
R9229 AVDD.n390 AVDD.n389 1.87264
R9230 AVDD.n1425 AVDD.n1421 1.87022
R9231 AVDD.n2524 AVDD.n2522 1.75943
R9232 AVDD.n1707 AVDD.n1315 1.71667
R9233 AVDD.n1427 AVDD.n1426 1.7131
R9234 AVDD.n1271 AVDD.n1264 1.70953
R9235 AVDD.n1296 AVDD.n1289 1.70953
R9236 AVDD.n1717 AVDD.n1715 1.70953
R9237 AVDD.n1481 AVDD.n1480 1.70953
R9238 AVDD.n3308 AVDD.n4 1.70953
R9239 AVDD.n1272 AVDD.n1248 1.70046
R9240 AVDD.n1297 AVDD.n1273 1.70046
R9241 AVDD.n1714 AVDD.n1713 1.70046
R9242 AVDD.n1708 AVDD.n1299 1.70046
R9243 AVDD.n1432 AVDD.n1298 1.70046
R9244 AVDD.n1486 AVDD.n0 1.70046
R9245 AVDD.n3309 AVDD.n2 1.70046
R9246 AVDD.n2630 AVDD.n1 1.70046
R9247 AVDD.t144 AVDD.n2165 1.63674
R9248 AVDD.n2353 AVDD.n2336 1.59407
R9249 AVDD.n1264 AVDD.n1249 1.54573
R9250 AVDD.n1289 AVDD.n1274 1.54573
R9251 AVDD.n1717 AVDD.n1716 1.54573
R9252 AVDD.n1480 AVDD.n1465 1.54573
R9253 AVDD.n4 AVDD.n3 1.54573
R9254 AVDD.n1426 AVDD.n1411 1.54216
R9255 AVDD.n1315 AVDD.n1300 1.53859
R9256 AVDD.n1425 AVDD.n1424 1.48486
R9257 AVDD.n1263 AVDD.n1262 1.48418
R9258 AVDD.n1288 AVDD.n1287 1.48418
R9259 AVDD.n1718 AVDD.n1246 1.48418
R9260 AVDD.n1314 AVDD.n1313 1.48418
R9261 AVDD.n1479 AVDD.n1478 1.48418
R9262 AVDD.n389 AVDD.n388 1.48418
R9263 AVDD.t8 AVDD.n2096 1.47311
R9264 AVDD.n1264 AVDD.n1263 1.42902
R9265 AVDD.n1289 AVDD.n1288 1.42902
R9266 AVDD.n1718 AVDD.n1717 1.42902
R9267 AVDD.n1480 AVDD.n1479 1.42902
R9268 AVDD.n389 AVDD.n4 1.42902
R9269 AVDD.n1315 AVDD.n1314 1.41979
R9270 AVDD.n1426 AVDD.n1425 1.41595
R9271 AVDD.n2754 AVDD.t15 1.30949
R9272 AVDD.n2576 AVDD.n2352 1.20764
R9273 AVDD.n2805 AVDD.t23 1.14587
R9274 AVDD.n1057 AVDD.n732 1.12991
R9275 AVDD.n1048 AVDD.n1047 1.12991
R9276 AVDD.t141 AVDD.n502 1.06405
R9277 AVDD.n1034 AVDD.t1 0.989054
R9278 AVDD.t35 AVDD.n2728 0.982243
R9279 AVDD.t18 AVDD.n2677 0.818619
R9280 AVDD.n214 AVDD.n212 0.753441
R9281 AVDD.n3089 AVDD.n3088 0.753441
R9282 AVDD.n3042 AVDD.n256 0.753441
R9283 AVDD.n3039 AVDD.n260 0.753441
R9284 AVDD.n305 AVDD.n302 0.753441
R9285 AVDD.n2988 AVDD.n2987 0.753441
R9286 AVDD.n2945 AVDD.n344 0.753441
R9287 AVDD.n2942 AVDD.n354 0.753441
R9288 AVDD.n408 AVDD.n406 0.753441
R9289 AVDD.n2896 AVDD.n2895 0.753441
R9290 AVDD.n2849 AVDD.n449 0.753441
R9291 AVDD.n2846 AVDD.n452 0.753441
R9292 AVDD.n1359 AVDD.n1358 0.753441
R9293 AVDD.n1363 AVDD.n1362 0.753441
R9294 AVDD.n1670 AVDD.n1669 0.753441
R9295 AVDD.n1666 AVDD.n1665 0.753441
R9296 AVDD.n1612 AVDD.n1447 0.753441
R9297 AVDD.n1609 AVDD.n1451 0.753441
R9298 AVDD.n1555 AVDD.n1498 0.753441
R9299 AVDD.n1552 AVDD.n1502 0.753441
R9300 AVDD.n2245 AVDD.n2244 0.753441
R9301 AVDD.n2253 AVDD.n2232 0.753441
R9302 AVDD.n2314 AVDD.n2313 0.753441
R9303 AVDD.n2318 AVDD.n2317 0.753441
R9304 AVDD.n2410 AVDD.n2409 0.753441
R9305 AVDD.n2401 AVDD.n2400 0.753441
R9306 AVDD.n2508 AVDD.n2458 0.753441
R9307 AVDD.n2463 AVDD.n2461 0.753441
R9308 AVDD.n2555 AVDD.n2554 0.753441
R9309 AVDD.n2559 AVDD.n2558 0.753441
R9310 AVDD.n2621 AVDD.n2620 0.753441
R9311 AVDD.n2625 AVDD.n2624 0.753441
R9312 AVDD.n1874 AVDD.n524 0.753441
R9313 AVDD.n1871 AVDD.n528 0.753441
R9314 AVDD.n1826 AVDD.n1825 0.753441
R9315 AVDD.n1160 AVDD.n1157 0.753441
R9316 AVDD.n1200 AVDD.n1198 0.753441
R9317 AVDD.n1776 AVDD.n1775 0.753441
R9318 AVDD.n2816 AVDD.n1949 0.753441
R9319 AVDD.n2404 AVDD.n2403 0.753441
R9320 AVDD.n2765 AVDD.n2013 0.753441
R9321 AVDD.n2465 AVDD.n2464 0.753441
R9322 AVDD.n2713 AVDD.n2082 0.753441
R9323 AVDD.n2709 AVDD.n2088 0.753441
R9324 AVDD.n2662 AVDD.n2151 0.753441
R9325 AVDD.n2658 AVDD.n2157 0.753441
R9326 AVDD.n3277 AVDD.n3276 0.753441
R9327 AVDD.n3273 AVDD.n3272 0.753441
R9328 AVDD.n3222 AVDD.n3221 0.753441
R9329 AVDD.n3218 AVDD.n3217 0.753441
R9330 AVDD.n3170 AVDD.n3169 0.753441
R9331 AVDD.n3166 AVDD.n3165 0.753441
R9332 AVDD.n933 AVDD.n932 0.753441
R9333 AVDD.n798 AVDD.n796 0.753441
R9334 AVDD.n877 AVDD.n833 0.753441
R9335 AVDD.n872 AVDD.n837 0.753441
R9336 AVDD.n615 AVDD.n568 0.753441
R9337 AVDD.n616 AVDD.n583 0.753441
R9338 AVDD.n660 AVDD.n573 0.753441
R9339 AVDD.n661 AVDD.n587 0.753441
R9340 AVDD.n1106 AVDD.n714 0.496226
R9341 AVDD.n2645 AVDD.t192 0.491372
R9342 AVDD.n1058 AVDD.n1056 0.376971
R9343 AVDD.n1049 AVDD.n745 0.376971
R9344 AVDD.n2690 AVDD.t29 0.327748
R9345 AVDD.n1106 AVDD.n713 0.324218
R9346 AVDD.n1714 AVDD.n1297 0.236753
R9347 AVDD.n1297 AVDD.n1272 0.236127
R9348 AVDD.n3309 AVDD.n1 0.236127
R9349 AVDD.n1298 AVDD.n0 0.214663
R9350 AVDD.n1272 AVDD 0.195393
R9351 AVDD.n1708 AVDD.n1298 0.17158
R9352 AVDD.n1714 AVDD.n1708 0.171267
R9353 AVDD AVDD.n3309 0.170327
R9354 AVDD.n1415 AVDD.n1414 0.16546
R9355 AVDD.n1253 AVDD.n1252 0.165423
R9356 AVDD.n1278 AVDD.n1277 0.165423
R9357 AVDD.n1725 AVDD.n1724 0.165423
R9358 AVDD.n1304 AVDD.n1303 0.165423
R9359 AVDD.n1469 AVDD.n1468 0.165423
R9360 AVDD.n395 AVDD.n382 0.165423
R9361 AVDD.n2741 AVDD.t32 0.164124
R9362 AVDD.n1841 AVDD.n1141 0.155087
R9363 AVDD.n1253 AVDD.n555 0.135601
R9364 AVDD.n1278 AVDD.n1196 0.135601
R9365 AVDD.n1726 AVDD.n1725 0.135601
R9366 AVDD.n1304 AVDD.n239 0.135601
R9367 AVDD.n1469 AVDD.n329 0.135601
R9368 AVDD.n396 AVDD.n395 0.135601
R9369 AVDD.n1415 AVDD.n279 0.135562
R9370 AVDD.n1256 AVDD.n1255 0.114786
R9371 AVDD.n1258 AVDD.n1256 0.114786
R9372 AVDD.n1254 AVDD.n1250 0.114786
R9373 AVDD.n1259 AVDD.n1250 0.114786
R9374 AVDD.n1269 AVDD.n1268 0.114786
R9375 AVDD.n1268 AVDD.n1267 0.114786
R9376 AVDD.n1281 AVDD.n1280 0.114786
R9377 AVDD.n1283 AVDD.n1281 0.114786
R9378 AVDD.n1279 AVDD.n1275 0.114786
R9379 AVDD.n1284 AVDD.n1275 0.114786
R9380 AVDD.n1294 AVDD.n1293 0.114786
R9381 AVDD.n1293 AVDD.n1292 0.114786
R9382 AVDD.n1722 AVDD.n1721 0.114786
R9383 AVDD.n1721 AVDD.n1720 0.114786
R9384 AVDD.n1723 AVDD.n1241 0.114786
R9385 AVDD.n1719 AVDD.n1241 0.114786
R9386 AVDD.n1711 AVDD.n1710 0.114786
R9387 AVDD.n1711 AVDD.n190 0.114786
R9388 AVDD.n1307 AVDD.n1306 0.114786
R9389 AVDD.n1309 AVDD.n1307 0.114786
R9390 AVDD.n1305 AVDD.n1301 0.114786
R9391 AVDD.n1310 AVDD.n1301 0.114786
R9392 AVDD.n1705 AVDD.n1704 0.114786
R9393 AVDD.n1704 AVDD.n1703 0.114786
R9394 AVDD.n1418 AVDD.n1417 0.114786
R9395 AVDD.n1420 AVDD.n1418 0.114786
R9396 AVDD.n1416 AVDD.n1412 0.114786
R9397 AVDD.n1421 AVDD.n1412 0.114786
R9398 AVDD.n1429 AVDD.n1410 0.114786
R9399 AVDD.n1433 AVDD.n1410 0.114786
R9400 AVDD.n1472 AVDD.n1471 0.114786
R9401 AVDD.n1474 AVDD.n1472 0.114786
R9402 AVDD.n1470 AVDD.n1466 0.114786
R9403 AVDD.n1475 AVDD.n1466 0.114786
R9404 AVDD.n1483 AVDD.n1464 0.114786
R9405 AVDD.n1487 AVDD.n1464 0.114786
R9406 AVDD.n393 AVDD.n392 0.114786
R9407 AVDD.n392 AVDD.n391 0.114786
R9408 AVDD.n394 AVDD.n383 0.114786
R9409 AVDD.n390 AVDD.n383 0.114786
R9410 AVDD.n3306 AVDD.n3305 0.114786
R9411 AVDD.n3305 AVDD.n3304 0.114786
R9412 AVDD.n2836 AVDD.n465 0.114786
R9413 AVDD.n2445 AVDD.n2368 0.114786
R9414 AVDD.n2522 AVDD.n2368 0.114786
R9415 AVDD.n2524 AVDD.n2523 0.114786
R9416 AVDD.n2523 AVDD.n2352 0.114786
R9417 AVDD.n2576 AVDD.n2575 0.114786
R9418 AVDD.n2575 AVDD.n2353 0.114786
R9419 AVDD.n1914 AVDD.t134 0.0823119
R9420 AVDD.n1270 AVDD.n1265 0.0805
R9421 AVDD.n1295 AVDD.n1290 0.0805
R9422 AVDD.n1712 AVDD.n1247 0.0805
R9423 AVDD.n1706 AVDD.n1316 0.0805
R9424 AVDD.n1431 AVDD.n1430 0.0805
R9425 AVDD.n1485 AVDD.n1484 0.0805
R9426 AVDD.n3307 AVDD.n5 0.0805
R9427 AVDD.n2629 AVDD.n2628 0.0805
R9428 AVDD.n1255 AVDD.n1251 0.0665714
R9429 AVDD.n1280 AVDD.n1276 0.0665714
R9430 AVDD.n1722 AVDD.n1242 0.0665714
R9431 AVDD.n1306 AVDD.n1302 0.0665714
R9432 AVDD.n1417 AVDD.n1413 0.0665714
R9433 AVDD.n1471 AVDD.n1467 0.0665714
R9434 AVDD.n393 AVDD.n384 0.0665714
R9435 AVDD AVDD.n0 0.0663
R9436 AVDD.n1258 AVDD.n1257 0.0522857
R9437 AVDD.n1269 AVDD.n1266 0.0522857
R9438 AVDD.n1283 AVDD.n1282 0.0522857
R9439 AVDD.n1294 AVDD.n1291 0.0522857
R9440 AVDD.n1720 AVDD.n1243 0.0522857
R9441 AVDD.n1710 AVDD.n1709 0.0522857
R9442 AVDD.n1309 AVDD.n1308 0.0522857
R9443 AVDD.n1705 AVDD.n1317 0.0522857
R9444 AVDD.n1420 AVDD.n1419 0.0522857
R9445 AVDD.n1429 AVDD.n1428 0.0522857
R9446 AVDD.n1474 AVDD.n1473 0.0522857
R9447 AVDD.n1483 AVDD.n1482 0.0522857
R9448 AVDD.n391 AVDD.n385 0.0522857
R9449 AVDD.n3306 AVDD.n6 0.0522857
R9450 AVDD.n1265 AVDD.n1248 0.0499324
R9451 AVDD.n1290 AVDD.n1273 0.0499324
R9452 AVDD.n1713 AVDD.n1712 0.0499324
R9453 AVDD.n1316 AVDD.n1299 0.0499324
R9454 AVDD.n1432 AVDD.n1431 0.0499324
R9455 AVDD.n1486 AVDD.n1485 0.0499324
R9456 AVDD.n5 AVDD.n2 0.0499324
R9457 AVDD.n2630 AVDD.n2629 0.0499324
R9458 AVDD.n982 AVDD.n773 0.0458461
R9459 AVDD.n957 AVDD.n781 0.0332381
R9460 AVDD.n1918 AVDD.n1895 0.0225877
R9461 AVDD.n1005 AVDD.n1004 0.0220827
R9462 AVDD.n1042 AVDD.n747 0.0220827
R9463 AVDD.n1089 AVDD.n1087 0.0220827
R9464 AVDD.n1107 AVDD.n712 0.0220827
R9465 AVDD.n2649 AVDD.n2173 0.0220517
R9466 AVDD.n968 AVDD.n782 0.0219797
R9467 AVDD.n943 AVDD.n789 0.0219797
R9468 AVDD.n935 AVDD.n934 0.0219797
R9469 AVDD.n921 AVDD.n803 0.0219797
R9470 AVDD.n913 AVDD.n803 0.0219797
R9471 AVDD.n913 AVDD.n912 0.0219797
R9472 AVDD.n902 AVDD.n816 0.0219797
R9473 AVDD.n894 AVDD.n893 0.0219797
R9474 AVDD.n885 AVDD.n884 0.0219797
R9475 AVDD.n884 AVDD.n830 0.0219797
R9476 AVDD.n873 AVDD.n836 0.0219797
R9477 AVDD.n863 AVDD.n862 0.0219797
R9478 AVDD.n854 AVDD.n848 0.0219797
R9479 AVDD.n995 AVDD.n993 0.0219286
R9480 AVDD.n995 AVDD.n994 0.0219286
R9481 AVDD.n1066 AVDD.n736 0.0219286
R9482 AVDD.n1099 AVDD.n1098 0.0219286
R9483 AVDD.n1104 AVDD.n1103 0.0219286
R9484 AVDD.n1012 AVDD.n1011 0.021783
R9485 AVDD.n1067 AVDD.n735 0.021631
R9486 AVDD.n1004 AVDD.n760 0.0214832
R9487 AVDD.n801 AVDD.n800 0.0213831
R9488 AVDD.n924 AVDD.n923 0.0213831
R9489 AVDD.n904 AVDD.n903 0.0210847
R9490 AVDD.n1926 AVDD.n483 0.0206243
R9491 AVDD.n1240 AVDD.n1239 0.0204607
R9492 AVDD.n2637 AVDD.n2188 0.020136
R9493 AVDD.n3126 AVDD.n3125 0.0199764
R9494 AVDD.n1937 AVDD.n1936 0.0192891
R9495 AVDD.n2826 AVDD.n2825 0.0192891
R9496 AVDD.n2811 AVDD.n1956 0.0192891
R9497 AVDD.n1988 AVDD.n1987 0.0192891
R9498 AVDD.n2002 AVDD.n2001 0.0192891
R9499 AVDD.n2776 AVDD.n2002 0.0192891
R9500 AVDD.n2760 AVDD.n2020 0.0192891
R9501 AVDD.n2046 AVDD.n2045 0.0192891
R9502 AVDD.n2722 AVDD.n2072 0.0192891
R9503 AVDD.n2710 AVDD.n2087 0.0192891
R9504 AVDD.n2101 AVDD.n2087 0.0192891
R9505 AVDD.n2119 AVDD.n2118 0.0192891
R9506 AVDD.n2671 AVDD.n2141 0.0192891
R9507 AVDD.n2659 AVDD.n2156 0.0192891
R9508 AVDD.n973 AVDD.n781 0.01925
R9509 AVDD.n1084 AVDD.n1083 0.0190851
R9510 AVDD.n1086 AVDD.n724 0.0190851
R9511 AVDD.n1938 AVDD.n1937 0.0190282
R9512 AVDD.n2775 AVDD.n2774 0.0190282
R9513 AVDD.n1074 AVDD.n1073 0.0189524
R9514 AVDD.n1071 AVDD.n717 0.0189524
R9515 AVDD.n1088 AVDD.n712 0.0187854
R9516 AVDD.n2789 AVDD.n1989 0.0187672
R9517 AVDD.n2788 AVDD.n2786 0.0187672
R9518 AVDD.n820 AVDD.n816 0.0186981
R9519 AVDD.n1103 AVDD.n715 0.0186548
R9520 AVDD.n2673 AVDD.n2672 0.0185063
R9521 AVDD.n834 AVDD.n830 0.0183998
R9522 AVDD.n876 AVDD.n875 0.0183998
R9523 AVDD.n2737 AVDD.n2047 0.0182453
R9524 AVDD.n2736 AVDD.n2734 0.0182453
R9525 AVDD.n812 AVDD.n807 0.0181014
R9526 AVDD.n904 AVDD.n815 0.0181014
R9527 AVDD.n2724 AVDD.n2723 0.0179843
R9528 AVDD.n800 AVDD.n795 0.0178031
R9529 AVDD.n2686 AVDD.n2120 0.0177234
R9530 AVDD.n2685 AVDD.n2683 0.0177234
R9531 AVDD.n972 AVDD.n968 0.0175048
R9532 AVDD.n2764 AVDD.n2763 0.0172015
R9533 AVDD.n2761 AVDD.n2019 0.0172015
R9534 AVDD.n2815 AVDD.n2814 0.0166795
R9535 AVDD.n2812 AVDD.n1955 0.0166795
R9536 AVDD.n1972 AVDD.n1971 0.0164186
R9537 AVDD.n1043 AVDD.n746 0.0160875
R9538 AVDD.n1046 AVDD.n1045 0.0160875
R9539 AVDD.n1055 AVDD.n1052 0.0159762
R9540 AVDD.n1054 AVDD.n734 0.0159762
R9541 AVDD.n2067 AVDD.n2066 0.0158967
R9542 AVDD.n992 AVDD.n991 0.0156786
R9543 AVDD.n1016 AVDD.n1015 0.015488
R9544 AVDD.n1013 AVDD.n1008 0.015488
R9545 AVDD.n935 AVDD.n794 0.0154165
R9546 AVDD.n1026 AVDD.n1025 0.015381
R9547 AVDD.n1029 AVDD.n1028 0.015381
R9548 AVDD.n2700 AVDD.n2102 0.0153747
R9549 AVDD.n2696 AVDD.n2104 0.0153747
R9550 AVDD.n2084 AVDD.n2083 0.0151138
R9551 AVDD.n2712 AVDD.n2086 0.0151138
R9552 AVDD.n2747 AVDD.n2034 0.0148528
R9553 AVDD.n2153 AVDD.n2152 0.0145919
R9554 AVDD.n2661 AVDD.n2155 0.0145919
R9555 AVDD.n2156 AVDD.n100 0.0145919
R9556 AVDD.n2798 AVDD.n1975 0.0143309
R9557 AVDD.n853 AVDD.n851 0.0142231
R9558 AVDD.n1950 AVDD.n1939 0.0140699
R9559 AVDD.n1953 AVDD.n1952 0.0140699
R9560 AVDD.n2393 AVDD.n2388 0.0139731
R9561 AVDD.n2415 AVDD.n2378 0.0139731
R9562 AVDD.n2435 AVDD.n2374 0.0139731
R9563 AVDD.n2503 AVDD.n2460 0.0139731
R9564 AVDD.n2489 AVDD.n2488 0.0139731
R9565 AVDD.n2549 AVDD.n2359 0.0139731
R9566 AVDD.n2561 AVDD.n2560 0.0139731
R9567 AVDD.n2561 AVDD.n2350 0.0139731
R9568 AVDD.n2587 AVDD.n2347 0.0139731
R9569 AVDD.n2615 AVDD.n2340 0.0139731
R9570 AVDD.n893 AVDD.n821 0.0139248
R9571 AVDD.n829 AVDD.n826 0.0139248
R9572 AVDD.n2515 AVDD.n2370 0.0137859
R9573 AVDD.n841 AVDD.n836 0.0136265
R9574 AVDD.n2438 AVDD.n2437 0.0135988
R9575 AVDD.n2443 AVDD.n2372 0.0135988
R9576 AVDD.n2014 AVDD.n2003 0.013548
R9577 AVDD.n2017 AVDD.n2016 0.013548
R9578 AVDD.n2606 AVDD.n2605 0.0134117
R9579 AVDD.n1016 AVDD.n1006 0.0133897
R9580 AVDD.n1025 AVDD.n753 0.0132976
R9581 AVDD.n2001 AVDD.n1990 0.0132871
R9582 AVDD.n2484 AVDD.n2483 0.0132246
R9583 AVDD.n2540 AVDD.n2539 0.0130374
R9584 AVDD.n862 AVDD.n842 0.0130298
R9585 AVDD.n2135 AVDD.n2134 0.0130261
R9586 AVDD.n2137 AVDD.n2133 0.0130261
R9587 AVDD.n971 AVDD.n969 0.013
R9588 AVDD.n991 AVDD.n767 0.013
R9589 AVDD.n2591 AVDD.n2588 0.0128503
R9590 AVDD.n2590 AVDD.n2343 0.0128503
R9591 AVDD.n1046 AVDD.n725 0.0127902
R9592 AVDD.n2061 AVDD.n2048 0.0127651
R9593 AVDD.n1070 AVDD.n734 0.0127024
R9594 AVDD.n2062 AVDD.n2061 0.0125042
R9595 AVDD.n2064 AVDD.n2060 0.0125042
R9596 AVDD.n2507 AVDD.n2506 0.012476
R9597 AVDD.n2504 AVDD.n2459 0.012476
R9598 AVDD.n526 AVDD.n525 0.0122801
R9599 AVDD.n1873 AVDD.n526 0.0122801
R9600 AVDD.n1873 AVDD.n1872 0.0122801
R9601 AVDD.n1864 AVDD.n534 0.0122801
R9602 AVDD.n1860 AVDD.n539 0.0122801
R9603 AVDD.n1852 AVDD.n539 0.0122801
R9604 AVDD.n1852 AVDD.n1851 0.0122801
R9605 AVDD.n1851 AVDD.n547 0.0122801
R9606 AVDD.n554 AVDD.n547 0.0122801
R9607 AVDD.n1840 AVDD.n1142 0.0122801
R9608 AVDD.n1149 AVDD.n1142 0.0122801
R9609 AVDD.n1831 AVDD.n1149 0.0122801
R9610 AVDD.n1827 AVDD.n1154 0.0122801
R9611 AVDD.n1816 AVDD.n1166 0.0122801
R9612 AVDD.n1816 AVDD.n1815 0.0122801
R9613 AVDD.n1815 AVDD.n1167 0.0122801
R9614 AVDD.n1806 AVDD.n1175 0.0122801
R9615 AVDD.n1802 AVDD.n1180 0.0122801
R9616 AVDD.n1794 AVDD.n1180 0.0122801
R9617 AVDD.n1794 AVDD.n1793 0.0122801
R9618 AVDD.n1793 AVDD.n1188 0.0122801
R9619 AVDD.n1195 AVDD.n1188 0.0122801
R9620 AVDD.n1784 AVDD.n1783 0.0122801
R9621 AVDD.n1783 AVDD.n1197 0.0122801
R9622 AVDD.n1774 AVDD.n1197 0.0122801
R9623 AVDD.n1774 AVDD.n1773 0.0122801
R9624 AVDD.n1764 AVDD.n1216 0.0122801
R9625 AVDD.n1762 AVDD.n1217 0.0122801
R9626 AVDD.n1224 AVDD.n1217 0.0122801
R9627 AVDD.n1753 AVDD.n1224 0.0122801
R9628 AVDD.n1751 AVDD.n1225 0.0122801
R9629 AVDD.n1742 AVDD.n1240 0.0122801
R9630 AVDD.n1742 AVDD.n1741 0.0122801
R9631 AVDD.n1741 AVDD.n1727 0.0122801
R9632 AVDD.n3107 AVDD.n195 0.0122801
R9633 AVDD.n3107 AVDD.n3106 0.0122801
R9634 AVDD.n3106 AVDD.n196 0.0122801
R9635 AVDD.n3097 AVDD.n3096 0.0122801
R9636 AVDD.n3087 AVDD.n217 0.0122801
R9637 AVDD.n3087 AVDD.n3086 0.0122801
R9638 AVDD.n3086 AVDD.n218 0.0122801
R9639 AVDD.n3077 AVDD.n226 0.0122801
R9640 AVDD.n3073 AVDD.n231 0.0122801
R9641 AVDD.n3065 AVDD.n3064 0.0122801
R9642 AVDD.n3064 AVDD.n240 0.0122801
R9643 AVDD.n247 AVDD.n240 0.0122801
R9644 AVDD.n258 AVDD.n257 0.0122801
R9645 AVDD.n3041 AVDD.n258 0.0122801
R9646 AVDD.n3041 AVDD.n3040 0.0122801
R9647 AVDD.n3032 AVDD.n266 0.0122801
R9648 AVDD.n3028 AVDD.n271 0.0122801
R9649 AVDD.n3020 AVDD.n3019 0.0122801
R9650 AVDD.n3019 AVDD.n280 0.0122801
R9651 AVDD.n287 AVDD.n280 0.0122801
R9652 AVDD.n300 AVDD.n299 0.0122801
R9653 AVDD.n2996 AVDD.n300 0.0122801
R9654 AVDD.n2996 AVDD.n2995 0.0122801
R9655 AVDD.n2986 AVDD.n308 0.0122801
R9656 AVDD.n2982 AVDD.n313 0.0122801
R9657 AVDD.n2974 AVDD.n313 0.0122801
R9658 AVDD.n2974 AVDD.n2973 0.0122801
R9659 AVDD.n2973 AVDD.n321 0.0122801
R9660 AVDD.n328 AVDD.n321 0.0122801
R9661 AVDD.n2964 AVDD.n2963 0.0122801
R9662 AVDD.n2963 AVDD.n330 0.0122801
R9663 AVDD.n337 AVDD.n330 0.0122801
R9664 AVDD.n2954 AVDD.n337 0.0122801
R9665 AVDD.n2954 AVDD.n2953 0.0122801
R9666 AVDD.n2944 AVDD.n2943 0.0122801
R9667 AVDD.n2943 AVDD.n353 0.0122801
R9668 AVDD.n2935 AVDD.n353 0.0122801
R9669 AVDD.n2933 AVDD.n360 0.0122801
R9670 AVDD.n2924 AVDD.n2923 0.0122801
R9671 AVDD.n2923 AVDD.n374 0.0122801
R9672 AVDD.n381 AVDD.n374 0.0122801
R9673 AVDD.n2914 AVDD.n381 0.0122801
R9674 AVDD.n2914 AVDD.n2913 0.0122801
R9675 AVDD.n404 AVDD.n403 0.0122801
R9676 AVDD.n2904 AVDD.n404 0.0122801
R9677 AVDD.n2904 AVDD.n2903 0.0122801
R9678 AVDD.n2903 AVDD.n405 0.0122801
R9679 AVDD.n2889 AVDD.n413 0.0122801
R9680 AVDD.n2880 AVDD.n421 0.0122801
R9681 AVDD.n2880 AVDD.n2879 0.0122801
R9682 AVDD.n2879 AVDD.n422 0.0122801
R9683 AVDD.n2870 AVDD.n430 0.0122801
R9684 AVDD.n2866 AVDD.n435 0.0122801
R9685 AVDD.n2858 AVDD.n435 0.0122801
R9686 AVDD.n2858 AVDD.n2857 0.0122801
R9687 AVDD.n2857 AVDD.n443 0.0122801
R9688 AVDD.n450 AVDD.n443 0.0122801
R9689 AVDD.n2848 AVDD.n450 0.0122801
R9690 AVDD.n2848 AVDD.n2847 0.0122801
R9691 AVDD.n2847 AVDD.n451 0.0122801
R9692 AVDD.n494 AVDD.n493 0.0122801
R9693 AVDD.n2134 AVDD.n2121 0.0122432
R9694 AVDD.n1831 AVDD.n1830 0.0121165
R9695 AVDD.n1828 AVDD.n1151 0.0121165
R9696 AVDD.n2412 AVDD.n2411 0.0121018
R9697 AVDD.n2414 AVDD.n2382 0.0121018
R9698 AVDD.n3283 AVDD.n3282 0.0119943
R9699 AVDD.n3282 AVDD.n109 0.0119943
R9700 AVDD.n3271 AVDD.n109 0.0119943
R9701 AVDD.n3269 AVDD.n111 0.0119943
R9702 AVDD.n3258 AVDD.n3257 0.0119943
R9703 AVDD.n3257 AVDD.n121 0.0119943
R9704 AVDD.n124 AVDD.n121 0.0119943
R9705 AVDD.n3246 AVDD.n124 0.0119943
R9706 AVDD.n3246 AVDD.n3245 0.0119943
R9707 AVDD.n3239 AVDD.n3238 0.0119943
R9708 AVDD.n3238 AVDD.n127 0.0119943
R9709 AVDD.n130 AVDD.n127 0.0119943
R9710 AVDD.n3227 AVDD.n130 0.0119943
R9711 AVDD.n3223 AVDD.n135 0.0119943
R9712 AVDD.n3211 AVDD.n143 0.0119943
R9713 AVDD.n3211 AVDD.n3210 0.0119943
R9714 AVDD.n3210 AVDD.n144 0.0119943
R9715 AVDD.n3199 AVDD.n148 0.0119943
R9716 AVDD.n3195 AVDD.n153 0.0119943
R9717 AVDD.n3188 AVDD.n153 0.0119943
R9718 AVDD.n3188 AVDD.n3187 0.0119943
R9719 AVDD.n3187 AVDD.n160 0.0119943
R9720 AVDD.n163 AVDD.n160 0.0119943
R9721 AVDD.n3176 AVDD.n3175 0.0119943
R9722 AVDD.n3175 AVDD.n165 0.0119943
R9723 AVDD.n3164 AVDD.n165 0.0119943
R9724 AVDD.n3164 AVDD.n3163 0.0119943
R9725 AVDD.n3152 AVDD.n170 0.0119943
R9726 AVDD.n3141 AVDD.n174 0.0119943
R9727 AVDD.n3141 AVDD.n3140 0.0119943
R9728 AVDD.n3140 AVDD.n175 0.0119943
R9729 AVDD.n3129 AVDD.n179 0.0119943
R9730 AVDD.n3125 AVDD.n184 0.0119943
R9731 AVDD.n189 AVDD.n184 0.0119943
R9732 AVDD.n3114 AVDD.n189 0.0119943
R9733 AVDD.n3112 AVDD.n191 0.0119943
R9734 AVDD.n1336 AVDD.n191 0.0119943
R9735 AVDD.n1344 AVDD.n1336 0.0119943
R9736 AVDD.n1355 AVDD.n1331 0.0119943
R9737 AVDD.n1357 AVDD.n1329 0.0119943
R9738 AVDD.n1368 AVDD.n1329 0.0119943
R9739 AVDD.n1370 AVDD.n1368 0.0119943
R9740 AVDD.n1381 AVDD.n1326 0.0119943
R9741 AVDD.n1385 AVDD.n1318 0.0119943
R9742 AVDD.n1701 AVDD.n1319 0.0119943
R9743 AVDD.n1694 AVDD.n1319 0.0119943
R9744 AVDD.n1694 AVDD.n1693 0.0119943
R9745 AVDD.n1676 AVDD.n1675 0.0119943
R9746 AVDD.n1675 AVDD.n1398 0.0119943
R9747 AVDD.n1664 AVDD.n1398 0.0119943
R9748 AVDD.n1662 AVDD.n1400 0.0119943
R9749 AVDD.n1651 AVDD.n1650 0.0119943
R9750 AVDD.n1644 AVDD.n1643 0.0119943
R9751 AVDD.n1643 AVDD.n1436 0.0119943
R9752 AVDD.n1439 AVDD.n1436 0.0119943
R9753 AVDD.n1621 AVDD.n1620 0.0119943
R9754 AVDD.n1620 AVDD.n1617 0.0119943
R9755 AVDD.n1617 AVDD.n1616 0.0119943
R9756 AVDD.n1611 AVDD.n1610 0.0119943
R9757 AVDD.n1603 AVDD.n1602 0.0119943
R9758 AVDD.n1602 AVDD.n1460 0.0119943
R9759 AVDD.n1463 AVDD.n1460 0.0119943
R9760 AVDD.n1591 AVDD.n1463 0.0119943
R9761 AVDD.n1591 AVDD.n1590 0.0119943
R9762 AVDD.n1584 AVDD.n1583 0.0119943
R9763 AVDD.n1583 AVDD.n1490 0.0119943
R9764 AVDD.n1493 AVDD.n1490 0.0119943
R9765 AVDD.n1572 AVDD.n1493 0.0119943
R9766 AVDD.n1572 AVDD.n1571 0.0119943
R9767 AVDD.n1554 AVDD.n1553 0.0119943
R9768 AVDD.n1553 AVDD.n1499 0.0119943
R9769 AVDD.n1546 AVDD.n1499 0.0119943
R9770 AVDD.n1544 AVDD.n1505 0.0119943
R9771 AVDD.n1533 AVDD.n1532 0.0119943
R9772 AVDD.n1532 AVDD.n1515 0.0119943
R9773 AVDD.n1520 AVDD.n1515 0.0119943
R9774 AVDD.n1521 AVDD.n1520 0.0119943
R9775 AVDD.n1521 AVDD.n7 0.0119943
R9776 AVDD.n3302 AVDD.n8 0.0119943
R9777 AVDD.n2236 AVDD.n8 0.0119943
R9778 AVDD.n2236 AVDD.n2233 0.0119943
R9779 AVDD.n2246 AVDD.n2233 0.0119943
R9780 AVDD.n2261 AVDD.n2258 0.0119943
R9781 AVDD.n2259 AVDD.n2228 0.0119943
R9782 AVDD.n2272 AVDD.n2228 0.0119943
R9783 AVDD.n2273 AVDD.n2272 0.0119943
R9784 AVDD.n2287 AVDD.n2279 0.0119943
R9785 AVDD.n2298 AVDD.n2223 0.0119943
R9786 AVDD.n2300 AVDD.n2298 0.0119943
R9787 AVDD.n2300 AVDD.n2299 0.0119943
R9788 AVDD.n2299 AVDD.n2220 0.0119943
R9789 AVDD.n2311 AVDD.n2220 0.0119943
R9790 AVDD.n2312 AVDD.n2311 0.0119943
R9791 AVDD.n2312 AVDD.n2218 0.0119943
R9792 AVDD.n2331 AVDD.n2218 0.0119943
R9793 AVDD.n2320 AVDD.n2215 0.0119943
R9794 AVDD.n1727 AVDD.n1726 0.0119529
R9795 AVDD.n2425 AVDD.n2424 0.0119147
R9796 AVDD.n1107 AVDD.n1106 0.0118909
R9797 AVDD.n787 AVDD.n782 0.0118365
R9798 AVDD.n946 AVDD.n945 0.0118365
R9799 AVDD.n3227 AVDD.n3226 0.0118346
R9800 AVDD.n3224 AVDD.n132 0.0118346
R9801 AVDD.n1106 AVDD.n1104 0.0118095
R9802 AVDD.n345 AVDD.n338 0.0117893
R9803 AVDD.n351 AVDD.n350 0.0117893
R9804 AVDD.n2626 AVDD.n2212 0.0117275
R9805 AVDD.n2018 AVDD.n2017 0.0117213
R9806 AVDD.n3114 AVDD.n3113 0.011675
R9807 AVDD.n2497 AVDD.n2472 0.0115404
R9808 AVDD.n1565 AVDD.n1494 0.0115153
R9809 AVDD.n1564 AVDD.n1560 0.0115153
R9810 AVDD.n3055 AVDD.n248 0.011462
R9811 AVDD.n3054 AVDD.n3050 0.011462
R9812 AVDD.n3005 AVDD.n290 0.011462
R9813 AVDD.n411 AVDD.n405 0.011462
R9814 AVDD.n2894 AVDD.n2893 0.011462
R9815 AVDD.n1773 AVDD.n1203 0.0112984
R9816 AVDD.n1215 AVDD.n1210 0.0112984
R9817 AVDD.n1954 AVDD.n1953 0.0111994
R9818 AVDD.n1687 AVDD.n1393 0.011196
R9819 AVDD.n1686 AVDD.n1682 0.011196
R9820 AVDD.n1627 AVDD.n1442 0.011196
R9821 AVDD.n2251 AVDD.n2246 0.011196
R9822 AVDD.n2252 AVDD.n2231 0.011196
R9823 AVDD.n2581 AVDD.n2580 0.0111662
R9824 AVDD.n1887 AVDD.n516 0.0111348
R9825 AVDD.n1886 AVDD.n1882 0.0111348
R9826 AVDD.n1784 AVDD.n1196 0.0111348
R9827 AVDD.n3163 AVDD.n167 0.0110364
R9828 AVDD.n3157 AVDD.n3156 0.0110364
R9829 AVDD.n2550 AVDD.n2358 0.010979
R9830 AVDD.n2553 AVDD.n2552 0.010979
R9831 AVDD.n3065 AVDD.n239 0.0109712
R9832 AVDD.n2801 AVDD.n1969 0.0109384
R9833 AVDD.n2800 AVDD.n2798 0.0109384
R9834 AVDD.n3291 AVDD.n102 0.0108768
R9835 AVDD.n3289 AVDD.n3288 0.0108768
R9836 AVDD.n3176 AVDD.n164 0.0108768
R9837 AVDD.n1895 AVDD.n477 0.0108076
R9838 AVDD.n1882 AVDD.n518 0.0108076
R9839 AVDD.n2493 AVDD.n2477 0.0107919
R9840 AVDD.n1702 AVDD.n1701 0.0107171
R9841 AVDD.n2661 AVDD.n2660 0.0106775
R9842 AVDD.n208 AVDD.n196 0.010644
R9843 AVDD.n210 AVDD.n204 0.010644
R9844 AVDD.n946 AVDD.n787 0.0106432
R9845 AVDD.n945 AVDD.n943 0.0106432
R9846 AVDD.n2616 AVDD.n2339 0.0106048
R9847 AVDD.n2619 AVDD.n2618 0.0106048
R9848 AVDD.n2173 AVDD.n100 0.0105575
R9849 AVDD.n3288 AVDD.n105 0.0105575
R9850 AVDD.n3050 AVDD.n250 0.0104804
R9851 AVDD.n3010 AVDD.n288 0.0104804
R9852 AVDD.n3009 AVDD.n3005 0.0104804
R9853 AVDD.n403 AVDD.n396 0.0104804
R9854 AVDD.n2429 AVDD.n2428 0.0104177
R9855 AVDD.n2750 AVDD.n2033 0.0104165
R9856 AVDD.n2749 AVDD.n2747 0.0104165
R9857 AVDD.n1344 AVDD.n1343 0.0103978
R9858 AVDD.n1341 AVDD.n1338 0.0103978
R9859 AVDD.n2995 AVDD.n301 0.0103167
R9860 AVDD.n1682 AVDD.n1396 0.0102382
R9861 AVDD.n1632 AVDD.n1440 0.0102382
R9862 AVDD.n1631 AVDD.n1627 0.0102382
R9863 AVDD.n3303 AVDD.n3302 0.0102382
R9864 AVDD.n2394 AVDD.n2385 0.0102305
R9865 AVDD.n2397 AVDD.n2396 0.0102305
R9866 AVDD.n2448 AVDD.n2447 0.0102305
R9867 AVDD.n2632 AVDD.n2631 0.0102305
R9868 AVDD.n2712 AVDD.n2711 0.0101555
R9869 AVDD.n352 AVDD.n351 0.0101531
R9870 AVDD.n1616 AVDD.n1445 0.0100785
R9871 AVDD.n2526 AVDD.n2525 0.0100434
R9872 AVDD.n1560 AVDD.n1497 0.0099189
R9873 AVDD.n2700 AVDD.n2699 0.00989457
R9874 AVDD.n2699 AVDD.n2103 0.00989457
R9875 AVDD.n2697 AVDD.n2103 0.00989457
R9876 AVDD.n2697 AVDD.n2696 0.00989457
R9877 AVDD.n2514 AVDD.n2454 0.00985629
R9878 AVDD.n2512 AVDD.n2511 0.00985629
R9879 AVDD.n1842 AVDD.n555 0.00982592
R9880 AVDD.n1083 AVDD.n725 0.00979257
R9881 AVDD.n1074 AVDD.n1070 0.00972619
R9882 AVDD.n1872 AVDD.n527 0.0096623
R9883 AVDD.n2711 AVDD.n2710 0.00963361
R9884 AVDD.n3239 AVDD.n125 0.00959962
R9885 AVDD.n1165 AVDD.n1154 0.00949869
R9886 AVDD.n458 AVDD.n451 0.00949869
R9887 AVDD.n2835 AVDD.n464 0.00948204
R9888 AVDD.n2601 AVDD.n2345 0.00948204
R9889 AVDD.n2597 AVDD.n2342 0.00948204
R9890 AVDD.n848 AVDD.n842 0.00944988
R9891 AVDD.n3271 AVDD.n3270 0.00943997
R9892 AVDD.n969 AVDD.n767 0.00942857
R9893 AVDD.n2066 AVDD.n2033 0.00937265
R9894 AVDD.n2750 AVDD.n2749 0.00937265
R9895 AVDD.n3040 AVDD.n259 0.00933508
R9896 AVDD.n2536 AVDD.n2535 0.00929491
R9897 AVDD.n142 AVDD.n135 0.00928033
R9898 AVDD.n2332 AVDD.n2331 0.00928033
R9899 AVDD.n1006 AVDD.n1005 0.00919305
R9900 AVDD.n2964 AVDD.n329 0.00917147
R9901 AVDD.n994 AVDD.n753 0.00913095
R9902 AVDD.n1664 AVDD.n1663 0.00912069
R9903 AVDD.n2660 AVDD.n2659 0.00911169
R9904 AVDD.n2531 AVDD.n2361 0.00910778
R9905 AVDD.n2935 AVDD.n2934 0.00900785
R9906 AVDD.n1584 AVDD.n1488 0.00896105
R9907 AVDD.n2602 AVDD.n2601 0.00892066
R9908 AVDD.n863 AVDD.n841 0.00885322
R9909 AVDD.n1971 AVDD.n1969 0.00885073
R9910 AVDD.n2801 AVDD.n2800 0.00885073
R9911 AVDD.n3020 AVDD.n279 0.00884424
R9912 AVDD.n420 AVDD.n413 0.00884424
R9913 AVDD.n1644 AVDD.n1434 0.00880141
R9914 AVDD.n1546 AVDD.n1545 0.00880141
R9915 AVDD.n2521 AVDD.n2369 0.00873353
R9916 AVDD.n1764 AVDD.n1763 0.00868063
R9917 AVDD.n2261 AVDD.n2260 0.00864176
R9918 AVDD.n2815 AVDD.n1954 0.00858977
R9919 AVDD.n826 AVDD.n821 0.00855489
R9920 AVDD.n885 AVDD.n829 0.00855489
R9921 AVDD.n2511 AVDD.n2455 0.00854641
R9922 AVDD.n3076 AVDD.n228 0.00851702
R9923 AVDD.n3074 AVDD.n3073 0.00851702
R9924 AVDD.n173 AVDD.n170 0.00848212
R9925 AVDD.n1174 AVDD.n1167 0.0083534
R9926 AVDD.n1382 AVDD.n1322 0.00832248
R9927 AVDD.n1385 AVDD.n1384 0.00832248
R9928 AVDD.n854 AVDD.n853 0.00825656
R9929 AVDD.n2397 AVDD.n2383 0.00817216
R9930 AVDD.n2530 AVDD.n2364 0.00817216
R9931 AVDD.n147 AVDD.n144 0.00816284
R9932 AVDD.n2764 AVDD.n2018 0.00806785
R9933 AVDD.n3096 AVDD.n211 0.00802618
R9934 AVDD.n2834 AVDD.n466 0.00798503
R9935 AVDD.n2420 AVDD.n2380 0.00798503
R9936 AVDD.n2429 AVDD.n2377 0.00798503
R9937 AVDD.n1237 AVDD.n1233 0.00786257
R9938 AVDD.n1356 AVDD.n1355 0.00784355
R9939 AVDD.n2577 AVDD.n2351 0.0077979
R9940 AVDD.n2619 AVDD.n2337 0.0077979
R9941 AVDD.n1841 AVDD.n1840 0.00769895
R9942 AVDD.n2986 AVDD.n2985 0.00769895
R9943 AVDD.n2983 AVDD.n310 0.00769895
R9944 AVDD.n429 AVDD.n422 0.00769895
R9945 AVDD.n2869 AVDD.n432 0.00769895
R9946 AVDD.n2867 AVDD.n2866 0.00769895
R9947 AVDD.n3128 AVDD.n181 0.00768391
R9948 AVDD.n2496 AVDD.n2473 0.00761078
R9949 AVDD.n2494 AVDD.n2493 0.00761078
R9950 AVDD.n1936 AVDD.n477 0.00754593
R9951 AVDD.n2683 AVDD.n2121 0.00754593
R9952 AVDD.n1753 AVDD.n1752 0.00753534
R9953 AVDD.n1610 AVDD.n1448 0.00752427
R9954 AVDD.n1459 AVDD.n1454 0.00752427
R9955 AVDD.n2273 AVDD.n2226 0.00752427
R9956 AVDD.n2286 AVDD.n2281 0.00752427
R9957 AVDD.n2284 AVDD.n2223 0.00752427
R9958 AVDD.n2446 AVDD.n2444 0.00742365
R9959 AVDD.n2553 AVDD.n2356 0.00742365
R9960 AVDD.n178 AVDD.n175 0.00736462
R9961 AVDD.n2062 AVDD.n2060 0.00728497
R9962 AVDD.n2724 AVDD.n2064 0.00728497
R9963 AVDD.n2573 AVDD.n2571 0.00723653
R9964 AVDD.n2581 AVDD.n2349 0.00723653
R9965 AVDD.n2838 AVDD.n463 0.00720811
R9966 AVDD.n1015 AVDD.n1008 0.00709472
R9967 AVDD.n1013 AVDD.n1012 0.00709472
R9968 AVDD.n794 AVDD.n789 0.00706325
R9969 AVDD.n2560 AVDD.n2356 0.0070494
R9970 AVDD.n1029 AVDD.n1026 0.00704762
R9971 AVDD.n1028 AVDD.n735 0.00704762
R9972 AVDD.n2335 AVDD.n2334 0.00704534
R9973 AVDD.n1864 AVDD.n1863 0.0070445
R9974 AVDD.n1861 AVDD.n536 0.0070445
R9975 AVDD.n1805 AVDD.n1177 0.0070445
R9976 AVDD.n1803 AVDD.n1802 0.0070445
R9977 AVDD.n2734 AVDD.n2048 0.00702401
R9978 AVDD.n118 AVDD.n111 0.0068857
R9979 AVDD.n120 AVDD.n114 0.0068857
R9980 AVDD.n3198 AVDD.n150 0.0068857
R9981 AVDD.n3196 AVDD.n3195 0.0068857
R9982 AVDD.n225 AVDD.n218 0.00688089
R9983 AVDD.n494 AVDD.n483 0.00688089
R9984 AVDD.n2497 AVDD.n2496 0.00686228
R9985 AVDD.n2494 AVDD.n2473 0.00686228
R9986 AVDD.n2135 AVDD.n2133 0.00676305
R9987 AVDD.n2673 AVDD.n2137 0.00676305
R9988 AVDD.n972 AVDD.n971 0.00675
R9989 AVDD.n993 AVDD.n992 0.00675
R9990 AVDD.n1370 AVDD.n1369 0.00672605
R9991 AVDD.n2320 AVDD.n2188 0.00672605
R9992 AVDD.n3032 AVDD.n3031 0.00671728
R9993 AVDD.n3029 AVDD.n268 0.00671728
R9994 AVDD.n1407 AVDD.n1400 0.00656641
R9995 AVDD.n1409 AVDD.n1403 0.00656641
R9996 AVDD.n2786 AVDD.n1990 0.00650209
R9997 AVDD.n1043 AVDD.n1042 0.0064952
R9998 AVDD.n1045 AVDD.n746 0.0064952
R9999 AVDD.n2424 AVDD.n2380 0.00648802
R10000 AVDD.n2420 AVDD.n2377 0.00648802
R10001 AVDD.n1052 AVDD.n736 0.00645238
R10002 AVDD.n1055 AVDD.n1054 0.00645238
R10003 AVDD.n371 AVDD.n360 0.00639005
R10004 AVDD.n371 AVDD.n367 0.00639005
R10005 AVDD.n373 AVDD.n367 0.00639005
R10006 AVDD.n2924 AVDD.n373 0.00639005
R10007 AVDD.n2387 AVDD.n466 0.0063009
R10008 AVDD.n2411 AVDD.n2383 0.0063009
R10009 AVDD.n1512 AVDD.n1505 0.00624713
R10010 AVDD.n1512 AVDD.n1508 0.00624713
R10011 AVDD.n1514 AVDD.n1508 0.00624713
R10012 AVDD.n1533 AVDD.n1514 0.00624713
R10013 AVDD.n2774 AVDD.n2003 0.00624113
R10014 AVDD.n2016 AVDD.n2014 0.00624113
R10015 AVDD.n3031 AVDD.n268 0.00606283
R10016 AVDD.n3029 AVDD.n3028 0.00606283
R10017 AVDD.n1407 AVDD.n1403 0.00592784
R10018 AVDD.n1651 AVDD.n1409 0.00592784
R10019 AVDD.n2507 AVDD.n2455 0.00592665
R10020 AVDD.n2627 AVDD.n2337 0.00592665
R10021 AVDD.n226 AVDD.n225 0.00589921
R10022 AVDD.n1369 AVDD.n1326 0.0057682
R10023 AVDD.n2521 AVDD.n2520 0.00573952
R10024 AVDD.n1863 AVDD.n536 0.0057356
R10025 AVDD.n1861 AVDD.n1860 0.0057356
R10026 AVDD.n1806 AVDD.n1805 0.0057356
R10027 AVDD.n1803 AVDD.n1177 0.0057356
R10028 AVDD.n2825 AVDD.n1939 0.00571921
R10029 AVDD.n1952 AVDD.n1950 0.00571921
R10030 AVDD.n118 AVDD.n114 0.00560856
R10031 AVDD.n3258 AVDD.n120 0.00560856
R10032 AVDD.n3199 AVDD.n3198 0.00560856
R10033 AVDD.n3196 AVDD.n150 0.00560856
R10034 AVDD.n2602 AVDD.n2343 0.0055524
R10035 AVDD.n1987 AVDD.n1975 0.00545825
R10036 AVDD.n2531 AVDD.n2530 0.00536527
R10037 AVDD.n2540 AVDD.n2361 0.00536527
R10038 AVDD.n1130 AVDD 0.00535819
R10039 AVDD.n1752 AVDD.n1751 0.00524476
R10040 AVDD.n2153 AVDD.n2141 0.00519729
R10041 AVDD.n2155 AVDD.n2152 0.00519729
R10042 AVDD.n2574 AVDD.n2351 0.00517814
R10043 AVDD.n179 AVDD.n178 0.00512963
R10044 AVDD.n1842 AVDD.n1841 0.00508115
R10045 AVDD.n2985 AVDD.n310 0.00508115
R10046 AVDD.n2983 AVDD.n2982 0.00508115
R10047 AVDD.n430 AVDD.n429 0.00508115
R10048 AVDD.n2870 AVDD.n2869 0.00508115
R10049 AVDD.n2867 AVDD.n432 0.00508115
R10050 AVDD.n2835 AVDD.n2834 0.00499102
R10051 AVDD.n2597 AVDD.n2345 0.00499102
R10052 AVDD.n2606 AVDD.n2342 0.00499102
R10053 AVDD.n1454 AVDD.n1448 0.00496999
R10054 AVDD.n1603 AVDD.n1459 0.00496999
R10055 AVDD.n2279 AVDD.n2226 0.00496999
R10056 AVDD.n2287 AVDD.n2286 0.00496999
R10057 AVDD.n2284 AVDD.n2281 0.00496999
R10058 AVDD.n2045 AVDD.n2034 0.00493633
R10059 AVDD.n1237 AVDD.n1225 0.00491754
R10060 AVDD.n1239 AVDD.n1233 0.00491754
R10061 AVDD.n3129 AVDD.n3128 0.00481034
R10062 AVDD.n3126 AVDD.n181 0.00481034
R10063 AVDD.n2444 AVDD.n2443 0.00480389
R10064 AVDD.n217 AVDD.n211 0.00475393
R10065 AVDD.n934 AVDD.n795 0.00467661
R10066 AVDD.n773 AVDD.n760 0.00467661
R10067 AVDD.n2084 AVDD.n2072 0.00467537
R10068 AVDD.n2086 AVDD.n2083 0.00467537
R10069 AVDD.n1357 AVDD.n1356 0.0046507
R10070 AVDD.n2515 AVDD.n2514 0.00461677
R10071 AVDD.n2512 AVDD.n2454 0.00461677
R10072 AVDD.n1175 AVDD.n1174 0.0044267
R10073 AVDD.n2102 AVDD.n2101 0.00441441
R10074 AVDD.n2118 AVDD.n2104 0.00441441
R10075 AVDD.n912 AVDD.n807 0.00437828
R10076 AVDD.n815 AVDD.n812 0.00437828
R10077 AVDD.n148 AVDD.n147 0.00433142
R10078 AVDD.n3077 AVDD.n3076 0.00426309
R10079 AVDD.n3074 AVDD.n228 0.00426309
R10080 AVDD.n2394 AVDD.n2393 0.00424252
R10081 AVDD.n2396 AVDD.n2385 0.00424252
R10082 AVDD.n2447 AVDD.n2369 0.00424252
R10083 AVDD.n1382 AVDD.n1381 0.00417178
R10084 AVDD.n1384 AVDD.n1322 0.00417178
R10085 AVDD.n1763 AVDD.n1762 0.00409948
R10086 AVDD.n876 AVDD.n834 0.00407995
R10087 AVDD.n875 AVDD.n873 0.00407995
R10088 AVDD.n851 AVDD.n760 0.00407995
R10089 AVDD.n1267 AVDD.n125 0.00407143
R10090 AVDD.n1292 AVDD.n164 0.00407143
R10091 AVDD.n3113 AVDD.n190 0.00407143
R10092 AVDD.n1703 AVDD.n1702 0.00407143
R10093 AVDD.n1434 AVDD.n1433 0.00407143
R10094 AVDD.n1488 AVDD.n1487 0.00407143
R10095 AVDD.n3304 AVDD.n3303 0.00407143
R10096 AVDD.n2428 AVDD.n2374 0.00405539
R10097 AVDD.n2354 AVDD.n2349 0.00405539
R10098 AVDD.n174 AVDD.n173 0.00401213
R10099 AVDD.n279 AVDD.n271 0.00393586
R10100 AVDD.n421 AVDD.n420 0.00393586
R10101 AVDD.n2067 AVDD.n2020 0.00389248
R10102 AVDD.n2578 AVDD.n2577 0.00386826
R10103 AVDD.n2616 AVDD.n2615 0.00386826
R10104 AVDD.n2618 AVDD.n2339 0.00386826
R10105 AVDD.n2260 AVDD.n2259 0.00385249
R10106 AVDD.n1089 AVDD.n1088 0.00379736
R10107 AVDD.n894 AVDD.n820 0.00378162
R10108 AVDD.n1099 AVDD.n715 0.00377381
R10109 AVDD.n2934 AVDD.n2933 0.00377225
R10110 AVDD.n1650 AVDD.n1434 0.00369285
R10111 AVDD.n1545 AVDD.n1544 0.00369285
R10112 AVDD.n2489 AVDD.n2477 0.00368114
R10113 AVDD.n2525 AVDD.n2367 0.00368114
R10114 AVDD.n2571 AVDD.n2354 0.00368114
R10115 AVDD.n1118 AVDD.n693 0.00365126
R10116 AVDD.n329 AVDD.n328 0.00360864
R10117 AVDD.n1590 AVDD.n1488 0.00353321
R10118 AVDD.n1084 AVDD.n724 0.0034976
R10119 AVDD.n1087 AVDD.n1086 0.0034976
R10120 AVDD.n2837 AVDD.n464 0.00349401
R10121 AVDD.n2550 AVDD.n2549 0.00349401
R10122 AVDD.n2552 AVDD.n2358 0.00349401
R10123 AVDD.n1073 AVDD.n1071 0.00347619
R10124 AVDD.n1098 AVDD.n717 0.00347619
R10125 AVDD.n266 AVDD.n259 0.00344503
R10126 AVDD.n1663 AVDD.n1662 0.00337356
R10127 AVDD.n1972 AVDD.n1956 0.00337056
R10128 AVDD.n2578 AVDD.n2350 0.00330689
R10129 AVDD.n2580 AVDD.n2347 0.00330689
R10130 AVDD.n1166 AVDD.n1165 0.00328141
R10131 AVDD.n2839 AVDD.n458 0.00328141
R10132 AVDD.n493 AVDD.n463 0.00328141
R10133 AVDD.n143 AVDD.n142 0.00321392
R10134 AVDD.n2332 AVDD.n2213 0.00321392
R10135 AVDD.n2334 AVDD.n2215 0.00321392
R10136 AVDD.n704 AVDD.n698 0.00321359
R10137 AVDD.n973 AVDD.n972 0.00317857
R10138 AVDD.n534 AVDD.n527 0.0031178
R10139 AVDD.n2814 AVDD.n1955 0.0031096
R10140 AVDD.n2812 AVDD.n2811 0.0031096
R10141 AVDD.n3270 AVDD.n3269 0.00305428
R10142 AVDD.n555 AVDD.n554 0.00295419
R10143 AVDD.n2472 AVDD.n2460 0.00293263
R10144 AVDD.n2526 AVDD.n2363 0.00293263
R10145 AVDD.n3245 AVDD.n125 0.00289464
R10146 AVDD.n2839 AVDD.n2838 0.00279058
R10147 AVDD.n2448 AVDD.n2446 0.00274551
R10148 AVDD.n2536 AVDD.n2363 0.00274551
R10149 AVDD.n2632 AVDD.n2212 0.00274551
R10150 AVDD.n2335 AVDD.n2213 0.00273499
R10151 AVDD.n2944 AVDD.n352 0.00262696
R10152 AVDD.n2763 AVDD.n2019 0.00258768
R10153 AVDD.n2761 AVDD.n2760 0.00258768
R10154 AVDD.n1554 AVDD.n1497 0.00257535
R10155 AVDD.n2838 AVDD.n2837 0.00255838
R10156 AVDD.n2425 AVDD.n2378 0.00255838
R10157 AVDD.n2574 AVDD.n2573 0.00255838
R10158 AVDD.n308 AVDD.n301 0.00246335
R10159 AVDD.n1611 AVDD.n1445 0.00241571
R10160 AVDD.n2412 AVDD.n2382 0.00237126
R10161 AVDD.n2415 AVDD.n2414 0.00237126
R10162 AVDD.n257 AVDD.n250 0.00229974
R10163 AVDD.n288 AVDD.n287 0.00229974
R10164 AVDD.n3010 AVDD.n3009 0.00229974
R10165 AVDD.n2913 AVDD.n396 0.00229974
R10166 AVDD.n1676 AVDD.n1396 0.00225607
R10167 AVDD.n1440 AVDD.n1439 0.00225607
R10168 AVDD.n1632 AVDD.n1631 0.00225607
R10169 AVDD.n3303 AVDD.n7 0.00225607
R10170 AVDD.n208 AVDD.n204 0.00213613
R10171 AVDD.n3097 AVDD.n210 0.00213613
R10172 AVDD.n1343 AVDD.n1338 0.00209642
R10173 AVDD.n1341 AVDD.n1331 0.00209642
R10174 AVDD.n2120 AVDD.n2119 0.00206576
R10175 AVDD.n2686 AVDD.n2685 0.00206576
R10176 AVDD.n2506 AVDD.n2459 0.00199701
R10177 AVDD.n2504 AVDD.n2503 0.00199701
R10178 AVDD.n515 AVDD.n477 0.00197251
R10179 AVDD.n525 AVDD.n518 0.00197251
R10180 AVDD.n3292 AVDD.n100 0.00193678
R10181 AVDD.n3283 AVDD.n105 0.00193678
R10182 AVDD.n702 AVDD.n684 0.00185679
R10183 AVDD.n1131 AVDD.n684 0.00185679
R10184 AVDD.n1131 AVDD.n1130 0.00185679
R10185 AVDD.n239 AVDD.n231 0.0018089
R10186 AVDD.n2723 AVDD.n2722 0.0018048
R10187 AVDD.n1702 AVDD.n1318 0.00177714
R10188 AVDD.n1271 AVDD.n1270 0.00175
R10189 AVDD.n1296 AVDD.n1295 0.00175
R10190 AVDD.n1715 AVDD.n1247 0.00175
R10191 AVDD.n1707 AVDD.n1706 0.00175
R10192 AVDD.n1430 AVDD.n1427 0.00175
R10193 AVDD.n1484 AVDD.n1481 0.00175
R10194 AVDD.n3308 AVDD.n3307 0.00175
R10195 AVDD.n2628 AVDD.n2336 0.00175
R10196 AVDD.n516 AVDD.n515 0.00164529
R10197 AVDD.n1887 AVDD.n1886 0.00164529
R10198 AVDD.n1196 AVDD.n1195 0.00164529
R10199 AVDD.n2588 AVDD.n2587 0.00162275
R10200 AVDD.n2591 AVDD.n2590 0.00162275
R10201 AVDD.n3292 AVDD.n3291 0.0016175
R10202 AVDD.n3289 AVDD.n102 0.0016175
R10203 AVDD.n164 AVDD.n163 0.0016175
R10204 AVDD.n2047 AVDD.n2046 0.00154384
R10205 AVDD.n2737 AVDD.n2736 0.00154384
R10206 AVDD.n1106 AVDD.n1105 0.00150665
R10207 AVDD.n1210 AVDD.n1203 0.00148168
R10208 AVDD.n1216 AVDD.n1215 0.00148168
R10209 AVDD.n3157 AVDD.n167 0.00145785
R10210 AVDD.n3156 AVDD.n3152 0.00145785
R10211 AVDD.n2535 AVDD.n2364 0.00143563
R10212 AVDD.n2539 AVDD.n2359 0.00143563
R10213 AVDD.n903 AVDD.n902 0.00139499
R10214 AVDD.n248 AVDD.n247 0.00131806
R10215 AVDD.n3055 AVDD.n3054 0.00131806
R10216 AVDD.n299 AVDD.n290 0.00131806
R10217 AVDD.n2894 AVDD.n411 0.00131806
R10218 AVDD.n2893 AVDD.n2889 0.00131806
R10219 AVDD.n1693 AVDD.n1393 0.00129821
R10220 AVDD.n1687 AVDD.n1686 0.00129821
R10221 AVDD.n1621 AVDD.n1442 0.00129821
R10222 AVDD.n2252 AVDD.n2251 0.00129821
R10223 AVDD.n2258 AVDD.n2231 0.00129821
R10224 AVDD.n2672 AVDD.n2671 0.00128288
R10225 AVDD.n2488 AVDD.n2483 0.0012485
R10226 AVDD.n2484 AVDD.n2367 0.0012485
R10227 AVDD.n2627 AVDD.n2626 0.0012485
R10228 AVDD.n924 AVDD.n801 0.00109666
R10229 AVDD.n923 AVDD.n921 0.00109666
R10230 AVDD.n2605 AVDD.n2340 0.00106138
R10231 AVDD.n1989 AVDD.n1988 0.00102192
R10232 AVDD.n2789 AVDD.n2788 0.00102192
R10233 AVDD.n2953 AVDD.n338 0.000990838
R10234 AVDD.n350 AVDD.n345 0.000990838
R10235 AVDD.n1105 AVDD.n693 0.000981443
R10236 AVDD.n1571 AVDD.n1494 0.000978927
R10237 AVDD.n1565 AVDD.n1564 0.000978927
R10238 AVDD.n1118 AVDD.n704 0.000937675
R10239 AVDD.n702 AVDD.n698 0.000937675
R10240 AVDD.n2437 AVDD.n2435 0.000874251
R10241 AVDD.n2438 AVDD.n2372 0.000874251
R10242 AVDD.n2631 AVDD.n2335 0.000874251
R10243 AVDD.n1726 AVDD.n195 0.000827225
R10244 AVDD.n3113 AVDD.n3112 0.000819285
R10245 AVDD.n1011 AVDD.n747 0.00079976
R10246 AVDD.n1067 AVDD.n1066 0.000797619
R10247 AVDD.n2826 AVDD.n1938 0.00076096
R10248 AVDD.n2776 AVDD.n2775 0.00076096
R10249 AVDD.n2388 AVDD.n2387 0.000687126
R10250 AVDD.n2520 AVDD.n2370 0.000687126
R10251 AVDD.n1141 AVDD 0.00067507
R10252 AVDD.n1830 AVDD.n1151 0.000663613
R10253 AVDD.n1828 AVDD.n1827 0.000663613
R10254 AVDD.n3226 AVDD.n132 0.000659642
R10255 AVDD.n3224 AVDD.n3223 0.000659642
R10256 VB3.n37 VB3.t17 235.565
R10257 VB3.n43 VB3.t28 235.565
R10258 VB3.n50 VB3.t29 235.565
R10259 VB3.n57 VB3.t1 235.565
R10260 VB3.n64 VB3.t13 235.565
R10261 VB3.n40 VB3.n39 208.996
R10262 VB3.n47 VB3.n46 208.996
R10263 VB3.n66 VB3.n35 208.994
R10264 VB3.n54 VB3.n52 208.994
R10265 VB3.n61 VB3.n59 208.994
R10266 VB3.n40 VB3.n38 205.859
R10267 VB3.n47 VB3.n45 205.859
R10268 VB3.n54 VB3.n53 205.857
R10269 VB3.n61 VB3.n60 205.857
R10270 VB3.n37 VB3.n36 205.238
R10271 VB3.n43 VB3.n42 205.238
R10272 VB3.n50 VB3.n49 205.238
R10273 VB3.n57 VB3.n56 205.238
R10274 VB3.n64 VB3.n63 205.238
R10275 VB3.n68 VB3.n67 204.857
R10276 VB3.n14 VB3.t35 114.392
R10277 VB3.n32 VB3.t37 103.459
R10278 VB3.n24 VB3.t39 103.459
R10279 VB3.n16 VB3.t38 103.459
R10280 VB3.n14 VB3.t36 87.566
R10281 VB3.n67 VB3.t6 28.5655
R10282 VB3.n67 VB3.t10 28.5655
R10283 VB3.n36 VB3.t24 28.5655
R10284 VB3.n36 VB3.t26 28.5655
R10285 VB3.n39 VB3.t2 28.5655
R10286 VB3.n39 VB3.t19 28.5655
R10287 VB3.n38 VB3.t8 28.5655
R10288 VB3.n38 VB3.t33 28.5655
R10289 VB3.n42 VB3.t4 28.5655
R10290 VB3.n42 VB3.t15 28.5655
R10291 VB3.n46 VB3.t12 28.5655
R10292 VB3.n46 VB3.t32 28.5655
R10293 VB3.n45 VB3.t31 28.5655
R10294 VB3.n45 VB3.t9 28.5655
R10295 VB3.n49 VB3.t21 28.5655
R10296 VB3.n49 VB3.t7 28.5655
R10297 VB3.n52 VB3.t14 28.5655
R10298 VB3.n52 VB3.t5 28.5655
R10299 VB3.n53 VB3.t27 28.5655
R10300 VB3.n53 VB3.t22 28.5655
R10301 VB3.n56 VB3.t20 28.5655
R10302 VB3.n56 VB3.t18 28.5655
R10303 VB3.n59 VB3.t0 28.5655
R10304 VB3.n59 VB3.t11 28.5655
R10305 VB3.n60 VB3.t16 28.5655
R10306 VB3.n60 VB3.t34 28.5655
R10307 VB3.n63 VB3.t30 28.5655
R10308 VB3.n63 VB3.t23 28.5655
R10309 VB3.n35 VB3.t3 28.5655
R10310 VB3.n35 VB3.t25 28.5655
R10311 VB3.n32 VB3.n31 21.9607
R10312 VB3.n33 VB3.n32 21.9607
R10313 VB3.n24 VB3.n23 21.9607
R10314 VB3.n25 VB3.n24 21.9607
R10315 VB3.n17 VB3.n16 21.9607
R10316 VB3.n16 VB3.n4 21.9607
R10317 VB3 VB3.n68 6.59201
R10318 VB3.n34 VB3.n33 4.50943
R10319 VB3.n15 VB3.n13 4.5005
R10320 VB3.n19 VB3.n18 4.5005
R10321 VB3.n21 VB3.n20 4.5005
R10322 VB3.n22 VB3.n3 4.5005
R10323 VB3.n27 VB3.n26 4.5005
R10324 VB3.n28 VB3.n2 4.5005
R10325 VB3.n30 VB3.n29 4.5005
R10326 VB3.n1 VB3.n0 4.5005
R10327 VB3.n7 VB3.n6 3.4105
R10328 VB3.n41 VB3.n37 2.18641
R10329 VB3.n44 VB3.n43 2.11889
R10330 VB3.n51 VB3.n50 2.11889
R10331 VB3.n58 VB3.n57 2.11889
R10332 VB3.n65 VB3.n64 2.11889
R10333 VB3.n13 VB3.n12 1.88261
R10334 VB3.n9 VB3.n8 1.71918
R10335 VB3.n8 VB3.n5 1.70602
R10336 VB3.n12 VB3.n11 1.70209
R10337 VB3.n10 VB3.n9 1.69771
R10338 VB3.n66 VB3.n65 1.26203
R10339 VB3.n62 VB3.n61 1.09471
R10340 VB3.n55 VB3.n54 1.09471
R10341 VB3.n48 VB3.n47 1.09471
R10342 VB3.n41 VB3.n40 1.09471
R10343 VB3.n68 VB3.n66 0.99936
R10344 VB3.n55 VB3.n51 0.534577
R10345 VB3.n15 VB3.n14 0.412155
R10346 VB3.n22 VB3.n21 0.2005
R10347 VB3.n30 VB3.n2 0.189786
R10348 VB3.n44 VB3.n41 0.168603
R10349 VB3.n51 VB3.n48 0.166567
R10350 VB3.n62 VB3 0.154973
R10351 VB3.n20 VB3.n3 0.132575
R10352 VB3.n29 VB3.n28 0.1255
R10353 VB3.n33 VB3.n1 0.105857
R10354 VB3.n18 VB3.n17 0.0987143
R10355 VB3.n31 VB3.n30 0.0915714
R10356 VB3.n21 VB3.n4 0.0844286
R10357 VB3.n19 VB3.n13 0.0759717
R10358 VB3.n20 VB3.n19 0.0759717
R10359 VB3.n27 VB3.n3 0.0759717
R10360 VB3.n28 VB3.n27 0.0759717
R10361 VB3.n29 VB3.n0 0.0759717
R10362 VB3.n34 VB3.n0 0.0759717
R10363 VB3.n58 VB3.n55 0.0688067
R10364 VB3.n65 VB3.n62 0.0688067
R10365 VB3.n48 VB3.n44 0.0680233
R10366 VB3.n26 VB3.n23 0.0665714
R10367 VB3.n26 VB3.n25 0.063
R10368 VB3.n25 VB3.n2 0.0522857
R10369 VB3.n23 VB3.n22 0.0487143
R10370 VB3.n18 VB3.n4 0.0308571
R10371 VB3 VB3.n34 0.0288019
R10372 VB3.n31 VB3.n1 0.0237143
R10373 VB3.n9 VB3.n7 0.0175856
R10374 VB3.n12 VB3.n5 0.0175856
R10375 VB3.n7 VB3.n5 0.0175856
R10376 VB3.n17 VB3.n15 0.0165714
R10377 VB3.n10 VB3 0.01366
R10378 VB3 VB3.n58 0.0133467
R10379 VB3.n11 VB3.n6 0.00881538
R10380 VB3.n8 VB3.n6 0.00881538
R10381 VB3.n11 VB3.n10 0.00881538
C0 VB2 a_4970_542# 0.00204f
C1 a_4970_n2468# AVDD 0.00396f
C2 AVDD a_4454_1009# 0.00716f
C3 AVDD a_1486_4980# 0.00588f
C4 VB2 a_4970_1638# 0.00204f
C5 VB3 a_3744_542# 0.00203f
C6 VB2 a_2712_4093# 0.00385f
C7 a_3744_n964# VB3 0.00588f
C8 a_10777_5531# a_10777_5228# 0.0205f
C9 VB3 a_3744_3472# 0.00588f
C10 a_11544_1111# VB2 0.144f
C11 VB3 a_1486_5597# 0.00666f
C12 AVDD a_3228_1638# 0.00418f
C13 a_10691_2488# VB2 0.0866f
C14 a_10691_2488# a_10691_1583# 0.0012f
C15 a_8985_205# VB4 0.0129f
C16 a_1486_n3085# VB1 0.00792f
C17 a_3744_n3085# VB2 0.00385f
C18 AVDD a_10519_5228# 0.0666f
C19 a_3228_n1581# VB2 0.00385f
C20 VB1 a_2002_3472# 0.00951f
C21 VB1 a_3744_6484# 0.00781f
C22 a_4454_n2468# VB3 0.00205f
C23 IREF a_8985_2488# 0.00505f
C24 VB3 a_4970_5597# 0.00775f
C25 a_2002_n3085# AVDD 0.00722f
C26 IREF a_9838_1583# 0.144f
C27 VB4 a_10777_6762# 0.145f
C28 a_1486_n1581# AVDD 0.00588f
C29 a_11544_2488# VB4 0.00487f
C30 a_2712_n2468# VB1 0.00938f
C31 AVDD a_1486_2724# 0.00981f
C32 a_2002_n964# AVDD 0.00513f
C33 VB3 a_2712_1638# 5.37e-19
C34 AVDD a_3228_5597# 0.00394f
C35 VB2 a_4454_4980# 0.00774f
C36 a_9828_n3072# a_10086_n3072# 0.0557f
C37 VB1 a_4970_2103# 0.0118f
C38 AVDD a_1486_542# 0.00852f
C39 AVDD a_2712_4980# 0.00385f
C40 VB1 a_8985_2488# 0.0165f
C41 AVDD a_3744_n77# 0.00648f
C42 VB2 a_3744_4093# 0.00385f
C43 a_4970_n964# VB3 0.00109f
C44 a_9838_1583# VB1 0.00302f
C45 VB2 a_1486_6484# 0.00666f
C46 VB1 a_2712_n77# 0.00932f
C47 VB3 a_4970_3472# 0.00109f
C48 AVDD a_4454_1638# 0.00418f
C49 VB3 a_2712_5597# 0.00334f
C50 AVDD a_2002_4093# 0.00515f
C51 a_3228_n964# VB1 0.00842f
C52 a_4970_n3085# VB2 0.00204f
C53 AVDD a_1486_4093# 0.00611f
C54 VB3 a_4454_542# 0.00205f
C55 a_4454_n1581# VB2 0.00108f
C56 VB1 a_3228_3472# 0.00857f
C57 VB1 a_4970_6484# 0.00727f
C58 VB2 a_4454_2724# 0.00108f
C59 VB3 a_4970_1009# 0.00109f
C60 IREF a_11544_1583# 0.144f
C61 a_3228_n3085# AVDD 0.00616f
C62 VB4 a_8132_2488# 0.00113f
C63 VB4 a_10777_6298# 0.151f
C64 a_9838_205# VB4 0.0686f
C65 a_2712_n1581# AVDD 0.00385f
C66 AVDD a_2712_2724# 0.00778f
C67 a_3744_n2468# VB1 0.00788f
C68 VB3 a_3744_1638# 0.00203f
C69 AVDD a_4454_5597# 0.00394f
C70 a_10519_6298# a_10777_6298# 0.0557f
C71 a_8132_1583# a_8132_2488# 0.0012f
C72 IREF a_11544_205# 3.01e-19
C73 AVDD a_4970_2724# 0.00778f
C74 VB1 a_2002_1638# 0.0166f
C75 AVDD a_3744_4980# 0.00385f
C76 a_2712_n3085# VB3 0.00334f
C77 VB2 a_4970_4093# 0.00204f
C78 a_2002_n1581# VB3 0.00666f
C79 VB2 a_2712_6484# 0.00281f
C80 VB3 a_3744_5597# 0.00483f
C81 AVDD a_1486_1009# 0.00922f
C82 AVDD a_3228_4093# 0.00408f
C83 a_4454_n964# VB1 0.00733f
C84 AVDD a_2002_542# 0.00756f
C85 AVDD a_4454_n77# 0.00648f
C86 VB1 a_4454_3472# 0.00748f
C87 a_1486_n2468# VB2 0.00666f
C88 a_11544_205# VB1 0.00114f
C89 VB1 a_2002_5597# 0.00937f
C90 VB1 a_3228_n77# 0.00836f
C91 VB3 a_3228_4980# 0.00492f
C92 a_4454_n3085# AVDD 0.00617f
C93 IREF a_8985_1111# 0.163f
C94 VB4 a_9838_2488# 0.00159f
C95 VB4 a_10777_5995# 0.151f
C96 a_3744_n1581# AVDD 0.00385f
C97 a_10691_1583# VB4 0.00302f
C98 VB2 VB4 2.51f
C99 a_4970_n2468# VB1 0.00733f
C100 AVDD a_3744_2724# 0.00778f
C101 VB3 a_4970_542# 0.00109f
C102 VB3 a_4970_1638# 0.00109f
C103 VB1 a_4454_1009# 0.0118f
C104 VB1 a_1486_4980# 0.00834f
C105 a_8985_1583# a_8985_2488# 0.0012f
C106 VB3 a_2712_4093# 0.00334f
C107 a_11544_2488# a_11544_1583# 0.0012f
C108 a_8132_1583# VB2 0.018f
C109 AVDD a_2002_2103# 0.00814f
C110 a_10691_205# VB4 0.0159f
C111 VB1 a_3228_1638# 0.0156f
C112 AVDD a_4970_4980# 0.00385f
C113 a_3744_n3085# VB3 0.00485f
C114 VB2 a_2002_3472# 0.00666f
C115 a_3228_n1581# VB3 0.00388f
C116 a_8985_1111# VB1 0.00374f
C117 VB2 a_3744_6484# 0.00281f
C118 VB3 a_3228_2724# 0.00107f
C119 AVDD a_2712_1009# 0.00716f
C120 a_2002_n3085# VB1 0.00888f
C121 AVDD a_4454_4093# 0.00408f
C122 a_1486_n1581# VB1 0.00834f
C123 AVDD VB1 0.104p
C124 AVDD a_2002_6484# 0.00555f
C125 VB1 a_1486_2724# 0.0152f
C126 a_2712_n2468# VB2 0.0028f
C127 a_2002_n964# VB1 0.00937f
C128 VB1 a_3228_5597# 0.00842f
C129 VB3 a_4454_4980# 0.00205f
C130 a_8985_1111# a_8985_205# 0.00119f
C131 IREF a_10691_1111# 0.159f
C132 VB4 a_10777_5531# 0.152f
C133 AVDD a_2712_542# 0.00649f
C134 a_4970_n1581# AVDD 0.00385f
C135 VB2 a_4970_2103# 0.00204f
C136 VB1 a_2712_4980# 0.00932f
C137 AVDD a_4970_n77# 0.00648f
C138 VB1 a_1486_542# 0.0157f
C139 a_10519_5995# a_10777_5995# 0.0557f
C140 VB2 a_8985_2488# 0.0866f
C141 a_9838_1583# a_9838_2488# 0.0012f
C142 VB1 a_3744_n77# 0.00781f
C143 VB3 a_3744_4093# 0.00483f
C144 a_8132_1583# a_8132_1111# 0.00931f
C145 a_9838_1583# VB2 0.0214f
C146 AVDD a_3228_2103# 0.00707f
C147 VB2 a_2712_n77# 0.00385f
C148 VB1 a_4454_1638# 0.0146f
C149 VB3 a_1486_n77# 0.00666f
C150 AVDD a_10777_6762# 0.0288f
C151 a_4970_n3085# VB3 0.00776f
C152 a_3228_n964# VB2 0.0028f
C153 VB1 a_2002_4093# 0.00937f
C154 VB1 a_1486_4093# 0.00841f
C155 a_4454_n1581# VB3 0.00872f
C156 VB2 a_3228_3472# 0.00281f
C157 VB2 a_4970_6484# 0.00871f
C158 VB3 a_4454_2724# 0.00205f
C159 a_3228_n3085# VB1 0.00794f
C160 a_2712_n1581# VB1 0.00932f
C161 AVDD a_1486_3472# 0.00697f
C162 VB3 a_2712_2103# 5.37e-19
C163 AVDD a_3228_6484# 0.00449f
C164 VB1 a_2712_2724# 0.0162f
C165 a_3744_n2468# VB2 0.0028f
C166 VB1 a_4454_5597# 0.00733f
C167 IREF a_8132_205# 0.00366f
C168 VB1 a_4970_2724# 0.0141f
C169 VB4 a_10777_5228# 0.152f
C170 a_2002_n2468# AVDD 0.00503f
C171 VB1 a_3744_4980# 0.00781f
C172 VB3 a_3228_1009# 0.00107f
C173 VB3 a_4970_4093# 0.00775f
C174 a_11544_1583# VB2 0.018f
C175 a_8985_1583# a_8985_1111# 0.00931f
C176 VB3 a_2712_6484# 0.00439f
C177 AVDD a_4454_2103# 0.00707f
C178 AVDD a_3228_542# 0.00649f
C179 VB1 a_1486_1009# 0.0129f
C180 AVDD a_10777_6298# 0.00735f
C181 VB1 a_2002_542# 0.0166f
C182 a_4454_n964# VB2 0.00774f
C183 AVDD a_3744_1009# 0.00716f
C184 VB1 a_3228_4093# 0.00842f
C185 a_9828_n3072# VB3 0.0941f
C186 VB1 a_4454_n77# 0.00727f
C187 VB2 a_4454_3472# 0.00774f
C188 a_8132_205# VB1 0.00114f
C189 a_11544_205# VB2 0.0908f
C190 VB2 a_3228_n77# 0.00385f
C191 a_2712_n964# AVDD 0.00406f
C192 a_4454_n3085# VB1 0.00685f
C193 VB3 a_2002_n77# 0.00666f
C194 AVDD a_2712_3472# 0.00494f
C195 a_3744_n1581# VB1 0.00781f
C196 VB3 a_3744_2103# 0.00203f
C197 AVDD a_4454_6484# 0.00451f
C198 VB1 a_3744_2724# 0.0147f
C199 VB2 a_4454_1009# 0.00108f
C200 VB2 a_1486_4980# 0.00666f
C201 a_4970_n2468# VB2 0.0087f
C202 IREF VB1 3.14f
C203 VB1 a_2002_2103# 0.0138f
C204 a_3228_n2468# AVDD 0.00396f
C205 a_11544_1111# VB4 0.00374f
C206 a_10691_2488# VB4 0.0599f
C207 VB1 a_4970_4980# 0.00727f
C208 a_1486_n3085# VB3 0.00666f
C209 a_10519_5531# a_10777_5531# 0.0557f
C210 a_9838_1583# a_9838_1111# 0.00931f
C211 a_8985_1111# VB2 0.00175f
C212 VB3 a_3744_6484# 0.00588f
C213 AVDD a_1486_1638# 0.0062f
C214 IREF a_8985_205# 0.0899f
C215 VB1 a_2712_1009# 0.0139f
C216 AVDD a_10777_5995# 0.00736f
C217 AVDD VB2 36.4f
C218 VB1 a_4454_4093# 0.00733f
C219 VB1 a_2002_6484# 0.0093f
C220 a_2712_n2468# VB3 0.00439f
C221 a_2002_n964# VB2 0.00666f
C222 IREF a_11544_2488# 0.0908f
C223 VB2 a_3228_5597# 0.00385f
C224 AVDD a_3744_542# 0.00649f
C225 a_9570_n3072# VB1 1.21e-21
C226 a_3744_n964# AVDD 0.00406f
C227 VB1 a_2712_542# 0.0167f
C228 a_4970_n1581# VB1 0.00727f
C229 AVDD a_3744_3472# 0.00494f
C230 VB3 a_4970_2103# 0.00109f
C231 AVDD a_1486_5597# 0.00597f
C232 VB1 a_4970_n77# 0.00727f
C233 VB2 a_2712_4980# 0.00281f
C234 a_8985_205# VB1 0.0606f
C235 VB2 a_3744_n77# 0.00385f
C236 VB1 a_3228_2103# 0.0129f
C237 a_4454_n2468# AVDD 0.00396f
C238 VB3 a_2712_n77# 0.00334f
C239 AVDD a_4970_5597# 0.00394f
C240 VB2 a_4454_1638# 0.00108f
C241 a_3228_n964# VB3 0.00492f
C242 a_11544_2488# VB1 0.0685f
C243 VB3 a_3228_3472# 0.00492f
C244 a_10691_1111# VB2 0.00509f
C245 a_10691_1583# a_10691_1111# 0.00931f
C246 AVDD a_2712_1638# 0.00418f
C247 VB3 a_4970_6484# 0.00109f
C248 a_3228_n3085# VB2 0.00385f
C249 AVDD a_10777_5531# 0.00737f
C250 a_2712_n1581# VB2 0.00385f
C251 VB1 a_1486_3472# 0.00856f
C252 VB1 a_3228_6484# 0.00836f
C253 a_3744_n2468# VB3 0.00588f
C254 a_10691_1111# a_10691_205# 0.00119f
C255 IREF a_8132_2488# 0.0908f
C256 IREF a_9838_205# 3.01e-19
C257 VB2 a_4454_5597# 0.00108f
C258 IREF a_8985_1583# 0.00511f
C259 VB4 a_10519_6762# 0.0898f
C260 a_4970_n964# AVDD 0.00406f
C261 VB2 a_4970_2724# 0.00204f
C262 a_2002_n2468# VB1 0.00937f
C263 AVDD a_4970_3472# 0.00494f
C264 a_1486_n964# AVDD 0.00609f
C265 AVDD a_2712_5597# 0.00394f
C266 a_10519_6762# a_10519_6298# 0.00305f
C267 VB2 a_3744_4980# 0.00281f
C268 AVDD a_4454_542# 0.00649f
C269 VB1 a_4454_2103# 0.0118f
C270 AVDD a_4970_1009# 0.00716f
C271 VB1 a_3228_542# 0.0157f
C272 AVDD a_2002_4980# 0.00492f
C273 VB1 a_8132_2488# 0.069f
C274 a_9838_205# VB1 0.00416f
C275 VB2 a_3228_4093# 0.00385f
C276 VB1 a_3744_1009# 0.0124f
C277 a_8985_1583# VB1 0.00374f
C278 a_4454_n964# VB3 0.00205f
C279 a_10519_5228# a_10777_5228# 0.0557f
C280 VB2 a_4454_n77# 0.00108f
C281 VB3 a_4454_3472# 0.00205f
C282 a_11544_1583# a_11544_1111# 0.00931f
C283 a_8132_205# VB2 0.0908f
C284 VB3 a_2002_5597# 0.00666f
C285 AVDD a_3744_1638# 0.00418f
C286 VB3 a_3228_n77# 0.00388f
C287 a_2712_n964# VB1 0.00938f
C288 a_4454_n3085# VB2 0.00108f
C289 AVDD a_10777_5228# 0.011f
C290 a_3744_n1581# VB2 0.00385f
C291 VB1 a_2712_3472# 0.00953f
C292 VB1 a_4454_6484# 0.00727f
C293 a_4970_n2468# VB3 0.00109f
C294 IREF a_9838_2488# 0.0908f
C295 a_11544_1111# a_11544_205# 0.00119f
C296 VB3 a_4454_1009# 0.00205f
C297 IREF a_10691_1583# 0.00174f
C298 IREF VB2 17.3f
C299 a_2712_n3085# AVDD 0.0062f
C300 VB4 a_10519_6298# 0.0931f
C301 a_2002_n1581# AVDD 0.00492f
C302 a_3228_n2468# VB1 0.00842f
C303 AVDD a_2002_2724# 0.00885f
C304 VB3 a_3228_1638# 0.00107f
C305 AVDD a_3744_5597# 0.00394f
C306 a_10777_6762# a_10777_6298# 0.00305f
C307 VB2 a_4970_4980# 0.00871f
C308 IREF a_10691_205# 0.0866f
C309 VB1 a_1486_1638# 0.0156f
C310 AVDD a_3228_4980# 0.00385f
C311 a_2002_n3085# VB3 0.00666f
C312 VB1 a_9838_2488# 0.0715f
C313 VB2 a_4454_4093# 0.00108f
C314 a_1486_n1581# VB3 0.00666f
C315 VB1 VB2 16.3f
C316 AVDD VB3 34.7f
C317 VB2 a_2002_6484# 0.00666f
C318 AVDD a_4970_542# 0.00649f
C319 a_8132_1111# a_8132_205# 0.00119f
C320 VB3 a_3228_5597# 0.00387f
C321 AVDD a_4970_1638# 0.00418f
C322 VB1 a_3744_542# 0.0151f
C323 AVDD a_2712_4093# 0.00408f
C324 a_3744_n964# VB1 0.00788f
C325 VB1 a_3744_3472# 0.00803f
C326 a_4970_n1581# VB2 0.00204f
C327 a_10691_205# VB1 0.0569f
C328 VB1 a_1486_5597# 0.00841f
C329 VB2 a_4970_n77# 0.00204f
C330 VB3 a_2712_4980# 0.00439f
C331 a_8985_205# VB2 0.00505f
C332 a_3744_n3085# AVDD 0.00616f
C333 IREF a_8132_1111# 0.0215f
C334 VB4 a_10519_5995# 0.093f
C335 VB3 a_3744_n77# 0.00485f
C336 VB4 a_8985_2488# 0.0569f
C337 a_3228_n1581# AVDD 0.00385f
C338 AVDD a_3228_2724# 0.00778f
C339 a_4454_n2468# VB1 0.00733f
C340 VB3 a_4454_1638# 0.00205f
C341 VB1 a_4970_5597# 0.00733f
C342 a_10519_6298# a_10519_5995# 0.0205f
C343 VB3 a_2002_4093# 0.00666f
C344 a_11544_2488# VB2 3.02e-19
C345 AVDD a_1486_2103# 0.00911f
C346 VB3 a_1486_4093# 0.00666f
C347 VB1 a_2712_1638# 0.0166f
C348 AVDD a_4454_4980# 0.00385f
C349 a_3228_n3085# VB3 0.00388f
C350 a_2712_n1581# VB3 0.00334f
C351 VB2 a_1486_3472# 0.00666f
C352 VB2 a_3228_6484# 0.00281f
C353 VB3 a_2712_2724# 5.37e-19
C354 AVDD a_2002_1009# 0.00824f
C355 VB3 a_4454_5597# 0.00871f
C356 AVDD a_3744_4093# 0.00408f
C357 a_4970_n964# VB1 0.00733f
C358 a_10086_n3072# VB2 5.57e-20
C359 VB3 a_4970_2724# 0.00109f
C360 AVDD a_1486_6484# 0.00658f
C361 VB1 a_4970_3472# 0.00748f
C362 a_1486_n964# VB1 0.00841f
C363 a_2002_n2468# VB2 0.00666f
C364 VB1 a_2712_5597# 0.00938f
C365 VB3 a_3744_4980# 0.00588f
C366 AVDD a_1486_n77# 0.00851f
C367 a_4970_n3085# AVDD 0.00615f
C368 IREF a_9838_1111# 0.0181f
C369 VB4 a_10519_5531# 0.0932f
C370 VB1 a_4454_542# 0.0146f
C371 a_4454_n1581# AVDD 0.00385f
C372 a_11544_1583# VB4 0.00374f
C373 VB2 a_4454_2103# 0.00108f
C374 AVDD a_4454_2724# 0.00778f
C375 VB1 a_2002_4980# 0.0093f
C376 VB1 a_4970_1009# 0.0118f
C377 a_10777_6298# a_10777_5995# 0.0205f
C378 VB2 a_8132_2488# 3.02e-19
C379 VB3 a_3228_4093# 0.00387f
C380 a_9838_205# VB2 0.0942f
C381 a_8985_1583# VB2 0.159f
C382 AVDD a_2712_2103# 0.00707f
C383 VB3 a_4454_n77# 0.00872f
C384 a_11544_205# VB4 0.0724f
C385 VB1 a_3744_1638# 0.0151f
C386 AVDD a_10519_6762# 0.0844f
C387 a_4454_n3085# VB3 0.00872f
C388 a_2712_n964# VB2 0.0028f
C389 a_3744_n1581# VB3 0.00485f
C390 VB2 a_2712_3472# 0.00281f
C391 a_9838_1111# VB1 0.00302f
C392 VB2 a_4454_6484# 0.00774f
C393 VB3 a_3744_2724# 0.00203f
C394 a_2712_n3085# VB1 0.0089f
C395 AVDD a_3228_1009# 0.00716f
C396 IREF VB3 0.00283f
C397 a_2002_n1581# VB1 0.0093f
C398 AVDD a_4970_4093# 0.00408f
C399 AVDD a_2712_6484# 0.00456f
C400 VB1 a_2002_2724# 0.0162f
C401 a_3228_n2468# VB2 0.0028f
C402 VB1 a_3744_5597# 0.00788f
C403 VB3 a_4970_4980# 0.00109f
C404 IREF a_11544_1111# 0.0181f
C405 IREF a_10691_2488# 0.00505f
C406 VB4 a_10519_5228# 0.0938f
C407 a_1486_n2468# AVDD 0.006f
C408 VB1 a_3228_4980# 0.00836f
C409 VB3 a_2712_1009# 5.37e-19
C410 a_10519_5995# a_10519_5531# 0.00305f
C411 VB2 a_9838_2488# 3.02e-19
C412 AVDD a_2002_n77# 0.00755f
C413 AVDD VB4 6.63f
C414 VB3 a_4454_4093# 0.00871f
C415 VB1 VB3 15.4f
C416 a_10691_1583# VB2 0.163f
C417 AVDD a_3744_2103# 0.00707f
C418 VB1 a_4970_542# 0.0146f
C419 VB1 a_4970_1638# 0.0146f
C420 AVDD a_10519_6298# 0.0631f
C421 VB1 a_2712_4093# 0.00938f
C422 a_9570_n3072# VB3 0.0941f
C423 a_3744_n964# VB2 0.0028f
C424 VB2 a_3744_3472# 0.00281f
C425 VB3 a_2712_542# 5.37e-19
C426 a_4970_n1581# VB3 0.00776f
C427 a_10691_205# VB2 0.00839f
C428 a_10691_2488# VB1 0.0132f
C429 VB3 a_4970_n77# 0.00776f
C430 a_3744_n3085# VB1 0.0074f
C431 a_1486_n3085# AVDD 0.00823f
C432 AVDD a_2002_3472# 0.00601f
C433 a_3228_n1581# VB1 0.00836f
C434 VB3 a_3228_2103# 0.00107f
C435 AVDD a_3744_6484# 0.00449f
C436 VB1 a_3228_2724# 0.0152f
C437 VB2 a_4970_5597# 0.00204f
C438 a_4454_n2468# VB2 0.00774f
C439 VB1 a_1486_2103# 0.0129f
C440 a_10691_1111# VB4 0.00302f
C441 a_2712_n2468# AVDD 0.00397f
C442 VB1 a_4454_4980# 0.00727f
C443 a_10777_5995# a_10777_5531# 0.00305f
C444 a_9838_1111# a_9838_205# 0.00119f
C445 a_8132_1111# VB2 0.144f
C446 AVDD a_4970_2103# 0.00707f
C447 VB3 a_3228_6484# 0.00492f
C448 VB1 a_2002_1009# 0.0139f
C449 AVDD a_10519_5995# 0.0631f
C450 a_4970_n964# VB2 0.0088f
C451 a_10086_n3072# VB3 0.15f
C452 VB1 a_3744_4093# 0.00788f
C453 VB1 a_1486_6484# 0.00834f
C454 VB2 a_4970_3472# 0.00871f
C455 AVDD a_2712_n77# 0.00648f
C456 a_1486_n964# VB2 0.00666f
C457 VB2 a_2712_5597# 0.00385f
C458 VB1 a_1486_n77# 0.00834f
C459 a_4970_n3085# VB1 0.00685f
C460 a_3228_n964# AVDD 0.00406f
C461 VB2 a_4454_542# 0.00108f
C462 AVDD a_3228_3472# 0.00494f
C463 a_4454_n1581# VB1 0.00727f
C464 VB3 a_4454_2103# 0.00205f
C465 AVDD a_4970_6484# 0.00448f
C466 VB1 a_4454_2724# 0.0141f
C467 VB3 a_3228_542# 0.00107f
C468 VB2 a_2002_4980# 0.00666f
C469 VB2 a_4970_1009# 0.00204f
C470 VB3 a_3744_1009# 0.00203f
C471 VB1 a_2712_2103# 0.0139f
C472 a_3744_n2468# AVDD 0.00396f
C473 a_8132_205# VB4 0.0686f
C474 a_2712_n964# VB3 0.00439f
C475 a_10519_5531# a_10519_5228# 0.0205f
C476 VB3 a_2712_3472# 0.00439f
C477 a_9838_1111# VB2 0.147f
C478 VB3 a_4454_6484# 0.00205f
C479 AVDD a_2002_1638# 0.00524f
C480 VB1 a_3228_1009# 0.0129f
C481 a_2712_n3085# VB2 0.00385f
C482 IREF VB4 1.36f
C483 AVDD a_10519_5531# 0.0631f
C484 VB1 a_4970_4093# 0.00733f
C485 VB1 a_2712_6484# 0.00932f
C486 a_3228_n2468# VB3 0.00492f
C487 IREF a_8132_1583# 0.147f
C488 VB2 a_3744_5597# 0.00385f
C489 a_4454_n964# AVDD 0.00406f
C490 a_1486_n2468# VB1 0.00841f
C491 AVDD a_4454_3472# 0.00494f
C492 AVDD a_2002_5597# 0.00501f
C493 a_10519_6762# a_10777_6762# 0.0557f
C494 VB2 a_3228_4980# 0.00281f
C495 AVDD a_3228_n77# 0.00648f
C496 a_9570_n3072# a_9828_n3072# 0.0557f
C497 VB1 a_2002_n77# 0.0093f
C498 VB2 VB3 27.5f
C499 VB1 VB4 4.15f
C500 VB1 a_3744_2103# 0.0123f
.ends

