** sch_path: /home/lci-ufsc/Desktop/work_sky130/INA_layout_v2/nfets_4x.sch
.subckt nfets_4x VS1 VS2 VB VG1 VG2 VD1 VD2
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
x1[2] VD1 VD2 VG2 VG1 VB VS2 VS1 nfets_2x
x1[1] VD1 VD2 VG2 VG1 VB VS2 VS1 nfets_2x
.ends

* expanding   symbol:  INA_layout_v2/nfets_2x.sym # of pins=7
** sym_path: /home/lci-ufsc/Desktop/work_sky130/INA_layout_v2/nfets_2x.sym
** sch_path: /home/lci-ufsc/Desktop/work_sky130/INA_layout_v2/nfets_2x.sch
.subckt nfets_2x VD1 VD2 VG2 VG1 VB VS2 VS1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
XM3[1] VB VB VB VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=9
XM3[0] VB VB VB VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=9
x1[2] VD1 VD2 VG2 VG1 VB VS2 VS1 nfets
x1[1] VD1 VD2 VG2 VG1 VB VS2 VS1 nfets
.ends


* expanding   symbol:  INA_layout_v2/nfets.sym # of pins=7
** sym_path: /home/lci-ufsc/Desktop/work_sky130/INA_layout_v2/nfets.sym
** sch_path: /home/lci-ufsc/Desktop/work_sky130/INA_layout_v2/nfets.sch
.subckt nfets VD1 VD2 VG2 VG1 VB VS2 VS1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
XM1 VD1 VG1 VS1 VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=7
XM2 VD2 VG2 VS2 VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=7
XM3 VB VB VB VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=4
.ends

.end
