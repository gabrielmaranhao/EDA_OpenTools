** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/ina_top.sch
.subckt ina_top IREF VI_1A VI_1B VI_2A VI_2B VO2 VO1 VCM AVDD AVSS
*.PININFO IREF:B VI_1A:B VI_1B:B VI_2A:B VI_2B:B VO2:B VO1:B VCM:B AVDD:B AVSS:B
x1 AVDD AVSS VI_1A VI_1B VO2 VO1 VCM VB1 VB2 VB3 VB4 VI_2A VI_2B dda
x2 IREF VB1 AVDD AVSS VB2 VB3 VB4 bias
.ends

* expanding   symbol:  INA_layout_v2/dda.sym # of pins=13
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/dda.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/dda.sch
.subckt dda AVDD AVSS VI_1A VI_1B VO2 VO1 VCM VB1 VB2 VB3 VB4 VI_2A VI_2B
*.PININFO AVDD:B VI_1A:B VI_1B:B VI_2A:B VI_2B:B VO1:B VO2:B VB1:B VB2:B VB3:B VB4:B VCM:B AVSS:B
x1 AVDD AVDD VB1 AVDD VB1 VIT_P2 VIT_P1 pfets_8x
x2 VIT_P1 VIT_P1 VI_1B AVDD VI_1A SUM_N SUM_P pfets_4x
x3 VIT_P2 VIT_P2 VI_2B AVDD VI_2A SUM_P SUM_N pfets_4x
x6 VD5 VD6 VB4 AVDD VB4 VO2 VO1 pfets_4x
x7 AVDD AVDD VCMFB AVDD VCMFB VD6 VD5 pfets_4x
x9 AVDD AVDD VD2 AVDD VD1 VD2 VD1 pfets_4x
x5 VO1 VO2 VB3 VB3 AVSS SUM_N SUM_P nfets_2x
x10 VD1 VCMFB VCM VO1 AVSS VIT_N1 VIT_N1 nfets_2x
x11 VD2 VCMFB VCM VO2 AVSS VIT_N2 VIT_N2 nfets_2x
x12 VIT_N1 VIT_N2 VB2 VB2 AVSS AVSS AVSS nfets_4x
x4 SUM_P SUM_N VB2 VB2 AVSS AVSS AVSS nfets_4x
x8 AVDD AVDD VCMFB AVDD VCMFB VCMFB VCMFB pfets_4x
.ends


* expanding   symbol:  INA_layout_v2/bias/bias.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/bias.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/bias.sch
.subckt bias IREF VB1 AVDD AVSS VB2 VB3 VB4
*.PININFO IREF:B VB1:B VB2:B VB3:B VB4:B AVDD:B AVSS:B
x1 IREF VB2 VB1 VB4 AVSS nbias_vb124
x2 VB3 VB1 VB2 AVDD pbias_vb123
x4 AVDD VB4 pbias_vb4
x3 VB3 AVSS nbias_vb3
.ends


* expanding   symbol:  INA_layout_v2/pfets_8x.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/pfets_8x.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/pfets_8x.sch
.subckt pfets_8x VS1 VS2 VG2 VB VG1 VD2 VD1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
x1[2] VS1 VS2 VG2 VB VG1 VD2 VD1 pfets_4x
x1[1] VS1 VS2 VG2 VB VG1 VD2 VD1 pfets_4x
.ends


* expanding   symbol:  INA_layout_v2/pfets_4x.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/pfets_4x.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/pfets_4x.sch
.subckt pfets_4x VS1 VS2 VG2 VB VG1 VD2 VD1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
x1[4] VS1 VS2 VG2 VB VG1 VD2 VD1 pfets
x1[3] VS1 VS2 VG2 VB VG1 VD2 VD1 pfets
x1[2] VS1 VS2 VG2 VB VG1 VD2 VD1 pfets
x1[1] VS1 VS2 VG2 VB VG1 VD2 VD1 pfets
.ends


* expanding   symbol:  INA_layout_v2/nfets_2x.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/nfets_2x.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/nfets_2x.sch
.subckt nfets_2x VD1 VD2 VG2 VG1 VB VS2 VS1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
XM3[1] VB VB VB VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=9
XM3[0] VB VB VB VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=9
x1[2] VD1 VD2 VG2 VG1 VB VS2 VS1 nfets
x1[1] VD1 VD2 VG2 VG1 VB VS2 VS1 nfets
.ends


* expanding   symbol:  INA_layout_v2/nfets_4x.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/nfets_4x.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/nfets_4x.sch
.subckt nfets_4x VD1 VD2 VG2 VG1 VB VS2 VS1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
x1[2] VD1 VD2 VG2 VG1 VB VS2 VS1 nfets_2x
x1[1] VD1 VD2 VG2 VG1 VB VS2 VS1 nfets_2x
.ends


* expanding   symbol:  INA_layout_v2/bias/nbias_vb124.sym # of pins=5
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/nbias_vb124.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/nbias_vb124.sch
.subckt nbias_vb124 IREF VB2 VB1 VB4 AVSS
*.PININFO IREF:B VB1:B VB2:B VB4:B AVSS:B
x1[5] AVSS AVSS IREF IREF nfet_2series
x1[4] AVSS AVSS IREF IREF nfet_2series
x1[3] AVSS AVSS IREF IREF nfet_2series
x1[2] AVSS AVSS IREF IREF nfet_2series
x1[1] AVSS AVSS IREF IREF nfet_2series
x2[5] AVSS AVSS IREF VB1 nfet_2series
x2[4] AVSS AVSS IREF VB1 nfet_2series
x2[3] AVSS AVSS IREF VB1 nfet_2series
x2[2] AVSS AVSS IREF VB1 nfet_2series
x2[1] AVSS AVSS IREF VB1 nfet_2series
x3[5] AVSS AVSS VB2 VB2 nfet_2series
x3[4] AVSS AVSS VB2 VB2 nfet_2series
x3[3] AVSS AVSS VB2 VB2 nfet_2series
x3[2] AVSS AVSS VB2 VB2 nfet_2series
x3[1] AVSS AVSS VB2 VB2 nfet_2series
x4[5] AVSS AVSS VB2 VB4 nfet_2series
x4[4] AVSS AVSS VB2 VB4 nfet_2series
x4[3] AVSS AVSS VB2 VB4 nfet_2series
x4[2] AVSS AVSS VB2 VB4 nfet_2series
x4[1] AVSS AVSS VB2 VB4 nfet_2series
XM1 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=44
.ends


* expanding   symbol:  INA_layout_v2/bias/pbias_vb123.sym # of pins=4
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/pbias_vb123.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/pbias_vb123.sch
.subckt pbias_vb123 VB3 VB1 VB2 AVDD
*.PININFO VB1:B VB2:B VB3:B AVDD:B
x1[35] AVDD AVDD VB1 VB1 pfet_2series
x1[34] AVDD AVDD VB1 VB1 pfet_2series
x1[33] AVDD AVDD VB1 VB1 pfet_2series
x1[32] AVDD AVDD VB1 VB1 pfet_2series
x1[31] AVDD AVDD VB1 VB1 pfet_2series
x1[30] AVDD AVDD VB1 VB1 pfet_2series
x1[29] AVDD AVDD VB1 VB1 pfet_2series
x1[28] AVDD AVDD VB1 VB1 pfet_2series
x1[27] AVDD AVDD VB1 VB1 pfet_2series
x1[26] AVDD AVDD VB1 VB1 pfet_2series
x1[25] AVDD AVDD VB1 VB1 pfet_2series
x1[24] AVDD AVDD VB1 VB1 pfet_2series
x1[23] AVDD AVDD VB1 VB1 pfet_2series
x1[22] AVDD AVDD VB1 VB1 pfet_2series
x1[21] AVDD AVDD VB1 VB1 pfet_2series
x1[20] AVDD AVDD VB1 VB1 pfet_2series
x1[19] AVDD AVDD VB1 VB1 pfet_2series
x1[18] AVDD AVDD VB1 VB1 pfet_2series
x1[17] AVDD AVDD VB1 VB1 pfet_2series
x1[16] AVDD AVDD VB1 VB1 pfet_2series
x1[15] AVDD AVDD VB1 VB1 pfet_2series
x1[14] AVDD AVDD VB1 VB1 pfet_2series
x1[13] AVDD AVDD VB1 VB1 pfet_2series
x1[12] AVDD AVDD VB1 VB1 pfet_2series
x1[11] AVDD AVDD VB1 VB1 pfet_2series
x1[10] AVDD AVDD VB1 VB1 pfet_2series
x1[9] AVDD AVDD VB1 VB1 pfet_2series
x1[8] AVDD AVDD VB1 VB1 pfet_2series
x1[7] AVDD AVDD VB1 VB1 pfet_2series
x1[6] AVDD AVDD VB1 VB1 pfet_2series
x1[5] AVDD AVDD VB1 VB1 pfet_2series
x1[4] AVDD AVDD VB1 VB1 pfet_2series
x1[3] AVDD AVDD VB1 VB1 pfet_2series
x1[2] AVDD AVDD VB1 VB1 pfet_2series
x1[1] AVDD AVDD VB1 VB1 pfet_2series
x2[35] AVDD AVDD VB1 VB3 pfet_2series
x2[34] AVDD AVDD VB1 VB3 pfet_2series
x2[33] AVDD AVDD VB1 VB3 pfet_2series
x2[32] AVDD AVDD VB1 VB3 pfet_2series
x2[31] AVDD AVDD VB1 VB3 pfet_2series
x2[30] AVDD AVDD VB1 VB3 pfet_2series
x2[29] AVDD AVDD VB1 VB3 pfet_2series
x2[28] AVDD AVDD VB1 VB3 pfet_2series
x2[27] AVDD AVDD VB1 VB3 pfet_2series
x2[26] AVDD AVDD VB1 VB3 pfet_2series
x2[25] AVDD AVDD VB1 VB3 pfet_2series
x2[24] AVDD AVDD VB1 VB3 pfet_2series
x2[23] AVDD AVDD VB1 VB3 pfet_2series
x2[22] AVDD AVDD VB1 VB3 pfet_2series
x2[21] AVDD AVDD VB1 VB3 pfet_2series
x2[20] AVDD AVDD VB1 VB3 pfet_2series
x2[19] AVDD AVDD VB1 VB3 pfet_2series
x2[18] AVDD AVDD VB1 VB3 pfet_2series
x2[17] AVDD AVDD VB1 VB3 pfet_2series
x2[16] AVDD AVDD VB1 VB3 pfet_2series
x2[15] AVDD AVDD VB1 VB3 pfet_2series
x2[14] AVDD AVDD VB1 VB3 pfet_2series
x2[13] AVDD AVDD VB1 VB3 pfet_2series
x2[12] AVDD AVDD VB1 VB3 pfet_2series
x2[11] AVDD AVDD VB1 VB3 pfet_2series
x2[10] AVDD AVDD VB1 VB3 pfet_2series
x2[9] AVDD AVDD VB1 VB3 pfet_2series
x2[8] AVDD AVDD VB1 VB3 pfet_2series
x2[7] AVDD AVDD VB1 VB3 pfet_2series
x2[6] AVDD AVDD VB1 VB3 pfet_2series
x2[5] AVDD AVDD VB1 VB3 pfet_2series
x2[4] AVDD AVDD VB1 VB3 pfet_2series
x2[3] AVDD AVDD VB1 VB3 pfet_2series
x2[2] AVDD AVDD VB1 VB3 pfet_2series
x2[1] AVDD AVDD VB1 VB3 pfet_2series
x3[35] AVDD AVDD VB1 VB2 pfet_2series
x3[34] AVDD AVDD VB1 VB2 pfet_2series
x3[33] AVDD AVDD VB1 VB2 pfet_2series
x3[32] AVDD AVDD VB1 VB2 pfet_2series
x3[31] AVDD AVDD VB1 VB2 pfet_2series
x3[30] AVDD AVDD VB1 VB2 pfet_2series
x3[29] AVDD AVDD VB1 VB2 pfet_2series
x3[28] AVDD AVDD VB1 VB2 pfet_2series
x3[27] AVDD AVDD VB1 VB2 pfet_2series
x3[26] AVDD AVDD VB1 VB2 pfet_2series
x3[25] AVDD AVDD VB1 VB2 pfet_2series
x3[24] AVDD AVDD VB1 VB2 pfet_2series
x3[23] AVDD AVDD VB1 VB2 pfet_2series
x3[22] AVDD AVDD VB1 VB2 pfet_2series
x3[21] AVDD AVDD VB1 VB2 pfet_2series
x3[20] AVDD AVDD VB1 VB2 pfet_2series
x3[19] AVDD AVDD VB1 VB2 pfet_2series
x3[18] AVDD AVDD VB1 VB2 pfet_2series
x3[17] AVDD AVDD VB1 VB2 pfet_2series
x3[16] AVDD AVDD VB1 VB2 pfet_2series
x3[15] AVDD AVDD VB1 VB2 pfet_2series
x3[14] AVDD AVDD VB1 VB2 pfet_2series
x3[13] AVDD AVDD VB1 VB2 pfet_2series
x3[12] AVDD AVDD VB1 VB2 pfet_2series
x3[11] AVDD AVDD VB1 VB2 pfet_2series
x3[10] AVDD AVDD VB1 VB2 pfet_2series
x3[9] AVDD AVDD VB1 VB2 pfet_2series
x3[8] AVDD AVDD VB1 VB2 pfet_2series
x3[7] AVDD AVDD VB1 VB2 pfet_2series
x3[6] AVDD AVDD VB1 VB2 pfet_2series
x3[5] AVDD AVDD VB1 VB2 pfet_2series
x3[4] AVDD AVDD VB1 VB2 pfet_2series
x3[3] AVDD AVDD VB1 VB2 pfet_2series
x3[2] AVDD AVDD VB1 VB2 pfet_2series
x3[1] AVDD AVDD VB1 VB2 pfet_2series
XM1 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=96
.ends


* expanding   symbol:  INA_layout_v2/bias/pbias_vb4.sym # of pins=2
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/pbias_vb4.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/pbias_vb4.sch
.subckt pbias_vb4 AVDD VB4
*.PININFO VB4:B AVDD:B
XM1 net1 VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM2 net2 VB4 net1 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM3 VB4 VB4 net2 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM4 net3 VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM5 net4 VB4 net3 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM6 VB4 VB4 net4 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM7 net5 VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM8 net6 VB4 net5 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM9 VB4 VB4 net6 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM10 net7 VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM11 net8 VB4 net7 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM12 VB4 VB4 net8 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM13 net9 VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM14 net10 VB4 net9 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM15 VB4 VB4 net10 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[20] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[19] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[18] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[17] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[16] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[15] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[14] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[13] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[12] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[11] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[10] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[9] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[8] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[7] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[6] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[5] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[4] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[3] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[2] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[1] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
.ends


* expanding   symbol:  INA_layout_v2/bias/nbias_vb3.sym # of pins=2
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/nbias_vb3.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/nbias_vb3.sch
.subckt nbias_vb3 VB3 AVSS
*.PININFO AVSS:B VB3:B
x1 AVSS AVSS VB3 net1 nfet_2series
x2 net1 AVSS VB3 VB3 nfet_2series
XM1[14] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[13] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[12] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[11] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[10] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[9] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[8] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[7] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[6] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[5] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[4] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[3] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[2] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[1] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
.ends


* expanding   symbol:  INA_layout_v2/pfets.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/pfets.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/pfets.sch
.subckt pfets VS1 VS2 VG2 VB VG1 VD2 VD1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
XM1 VD1 VG1 VS1 VB sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=22
XM2 VD2 VG2 VS2 VB sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=22
XM3 VB VB VB VB sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=34
.ends


* expanding   symbol:  INA_layout_v2/nfets.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/nfets.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/nfets.sch
.subckt nfets VD1 VD2 VG2 VG1 VB VS2 VS1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
XM1 VD1 VG1 VS1 VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=7
XM2 VD2 VG2 VS2 VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=7
XM3 VB VB VB VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=4
.ends


* expanding   symbol:  INA_layout_v2/bias/nfet_2series.sym # of pins=4
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/nfet_2series.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/nfet_2series.sch
.subckt nfet_2series S B G D
*.PININFO S:B B:B G:B D:B
XM1 D G net1 B sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM2 net1 G S B sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
.ends


* expanding   symbol:  INA_layout_v2/bias/pfet_2series.sym # of pins=4
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/pfet_2series.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/pfet_2series.sch
.subckt pfet_2series S B G D
*.PININFO S:B B:B G:B D:B
XM1 net1 G S B sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM2 D G net1 B sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
.ends

.end
