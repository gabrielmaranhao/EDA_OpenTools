** sch_path: /home/gmaranhao/pdk/IHP-Open-PDK/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/dc_lv_nmos.sch
**.subckt dc_lv_nmos
Vgs net1 GND 0.75
Vds net3 GND 1.5
XM1 net2 net1 GND GND sg13_lv_nmos W=1.0u L=0.45u ng=1 m=1
Vd net3 net2 0
.save i(vd)
**** begin user architecture code
 .lib /home/gmaranhao/pdk/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt



.param temp=27
.control
pre_osdi ./psp103_nqs.osdi
save all
op
*reset
dc Vds 0 3 0.01 Vgs 0. 0.9 0.1
write dc_lv_nmos.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
