** sch_path: /home/gmaranhao/Desktop/ihp130_work/PSPvsACM.sch
**.subckt PSPvsACM
VG vg GND 0
VD1 vd GND {vd}
VB net1 GND 0
VS net2 GND 0
N1 net4 vg net5 net3 NMOS_ACM w=10u l=0.12u n=1.414 is=11.77u vt0=0.4902 sigma=53.4m zeta=7m
VB3 net3 GND 0
VS_acm net5 GND 0
VD2 net4 GND {vd}
XM1 vd vg net2 net1 sg13_lv_nmos W=10.0u L=0.12u ng=1 m=1
**** begin user architecture code



.param vd=1.5

.control
pre_osdi ./psp103_nqs.osdi
pre_osdi /home/gmaranhao/Desktop/gf180_work/ACM/NMOS_ACM_2V0.osdi
save all



dc VG 0 1.5 1m
*let gm = deriv(i(vs))
*save gm
remzerovec
write PSPvsACM.raw
set appendwrite

*dc VG1 0 1.5 10m
*let gm = deriv(i(vs_acm))
*save gm
*remzerovec
*write PSPvsACM.raw

.endc



.lib /home/gmaranhao/pdk/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.model NMOS_ACM nmos_ACM

**** end user architecture code
**.ends
.GLOBAL GND
.end
